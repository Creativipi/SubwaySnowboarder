----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08.06.2025 00:00:57
-- Design Name: 
-- Module Name: BackMgmt - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity BackMgmt is
    Port ( 
        i_view_x : in STD_LOGIC_VECTOR (9 downto 0); -- position x du pixel � voir
        i_view_y : in STD_LOGIC_VECTOR (9 downto 0); -- position y du pixel � voir
        i_ch_we_tileBack : in STD_LOGIC;
        i_col : in STD_LOGIC_VECTOR (6 downto 0); -- prochaine tuile � changer
        i_row : in STD_LOGIC_VECTOR (6 downto 0); -- prochaine tuile � changer
        i_tile_id : in STD_LOGIC_VECTOR (4 downto 0); -- tuile qui change
        i_flip_y : in STD_LOGIC; -- valeur du flip
        i_ch_tile_id : in STD_LOGIC; -- change la tuile?
        i_ch_flipY : in STD_LOGIC; -- change le flip?
        i_clk : in STD_LOGIC; -- la clock

        -- Info du pixel qu'on regarde
        o_tile_id : out STD_LOGIC_VECTOR (4 downto 0); 
        o_flip_y : out STD_LOGIC;
        o_pix_x : out STD_LOGIC_VECTOR (2 downto 0);
        o_pix_y : out STD_LOGIC_VECTOR (2 downto 0)
    );
end BackMgmt;

architecture Behavioral of BackMgmt is

    signal s_view_index : std_logic_vector (13 downto 0);
    signal r_view_x, r_view_y : std_logic_vector(9 downto 0);

    -- Packed format: [5] = flip_y, [4:0] = tile_id
    type tile_data_array_t is array (0 to 16383) of std_logic_vector(5 downto 0);
    signal tile_data_map : tile_data_array_t := (
        1 => "000010",
129 => "000010",
257 => "000010",
385 => "000010",
513 => "000010",
641 => "000010",
769 => "000010",
897 => "000010",
1025 => "000010",
1153 => "000010",
1281 => "000010",
1409 => "000010",
1537 => "000010",
1665 => "000010",
1793 => "000010",
1921 => "000010",
2049 => "000010",
2177 => "000010",
2305 => "000010",
2433 => "000010",
2561 => "000010",
2689 => "000010",
2817 => "000010",
2945 => "000010",
3073 => "000010",
3201 => "000010",
3329 => "000010",
3457 => "000010",
3585 => "000010",
3713 => "000010",
3841 => "000010",
3969 => "000010",
4097 => "000010",
4225 => "000010",
4353 => "000010",
4481 => "000010",
4609 => "000010",
4737 => "000010",
4865 => "000010",
4993 => "000010",
5121 => "000010",
5249 => "000010",
5377 => "000010",
5505 => "000010",
5633 => "000010",
5761 => "000010",
5889 => "000010",
6017 => "000010",
6145 => "000010",
6273 => "000010",
6401 => "000010",
6529 => "000010",
6657 => "000010",
6785 => "000010",
6913 => "000010",
7041 => "000010",
7169 => "000010",
7297 => "000010",
7425 => "000010",
7553 => "000010",
7681 => "000010",
7809 => "000010",
7937 => "000010",
8065 => "000010",
8193 => "000010",
8321 => "000010",
8449 => "000010",
8577 => "000010",
8705 => "000010",
8833 => "000010",
8961 => "000010",
9089 => "000010",
9217 => "000010",
9345 => "000010",
9473 => "000010",
9601 => "000010",
9729 => "000010",
9857 => "000010",
9985 => "000010",
10113 => "000010",
10241 => "000010",
10369 => "000010",
10497 => "000010",
10625 => "000010",
10753 => "000010",
10881 => "000010",
11009 => "000010",
11137 => "000010",
11265 => "000010",
11393 => "000010",
11521 => "000010",
11649 => "000010",
11777 => "000010",
11905 => "000010",
12033 => "000010",
12161 => "000010",
12289 => "000010",
12417 => "000010",
12545 => "000010",
12673 => "000010",
12801 => "000010",
12929 => "000010",
13057 => "000010",
13185 => "000010",
13313 => "000010",
13441 => "000010",
13569 => "000010",
13697 => "000010",
13825 => "000010",
13953 => "000010",
14081 => "000010",
14209 => "000010",
14337 => "000010",
14465 => "000010",
14593 => "000010",
14721 => "000010",
14849 => "000010",
14977 => "000010",
15105 => "000010",
15233 => "000010",
15361 => "000010",
15489 => "000010",
15617 => "000010",
15745 => "000010",
15873 => "000010",
16001 => "000010",
16129 => "000010",
16257 => "000010",
7 => "000001",
135 => "000001",
263 => "000001",
391 => "000001",
519 => "000001",
647 => "000001",
775 => "000001",
903 => "000001",
1031 => "000001",
1159 => "000001",
1287 => "000001",
1415 => "000001",
1543 => "000001",
1671 => "000001",
1799 => "000001",
1927 => "000001",
2055 => "000001",
2183 => "000001",
2311 => "000001",
2439 => "000001",
2567 => "000001",
2695 => "000001",
2823 => "000001",
2951 => "000001",
3079 => "000001",
3207 => "000001",
3335 => "000001",
3463 => "000001",
3591 => "000001",
3719 => "000001",
3847 => "000001",
3975 => "000001",
4103 => "000001",
4231 => "000001",
4359 => "000001",
4487 => "000001",
4615 => "000001",
4743 => "000001",
4871 => "000001",
4999 => "000001",
5127 => "000001",
5255 => "000001",
5383 => "000001",
5511 => "000001",
5639 => "000001",
5767 => "000001",
5895 => "000001",
6023 => "000001",
6151 => "000001",
6279 => "000001",
6407 => "000001",
6535 => "000001",
6663 => "000001",
6791 => "000001",
6919 => "000001",
7047 => "000001",
7175 => "000001",
7303 => "000001",
7431 => "000001",
7559 => "000001",
7687 => "000001",
7815 => "000001",
7943 => "000001",
8071 => "000001",
8199 => "000001",
8327 => "000001",
8455 => "000001",
8583 => "000001",
8711 => "000001",
8839 => "000001",
8967 => "000001",
9095 => "000001",
9223 => "000001",
9351 => "000001",
9479 => "000001",
9607 => "000001",
9735 => "000001",
9863 => "000001",
9991 => "000001",
10119 => "000001",
10247 => "000001",
10375 => "000001",
10503 => "000001",
10631 => "000001",
10759 => "000001",
10887 => "000001",
11015 => "000001",
11143 => "000001",
11271 => "000001",
11399 => "000001",
11527 => "000001",
11655 => "000001",
11783 => "000001",
11911 => "000001",
12039 => "000001",
12167 => "000001",
12295 => "000001",
12423 => "000001",
12551 => "000001",
12679 => "000001",
12807 => "000001",
12935 => "000001",
13063 => "000001",
13191 => "000001",
13319 => "000001",
13447 => "000001",
13575 => "000001",
13703 => "000001",
13831 => "000001",
13959 => "000001",
14087 => "000001",
14215 => "000001",
14343 => "000001",
14471 => "000001",
14599 => "000001",
14727 => "000001",
14855 => "000001",
14983 => "000001",
15111 => "000001",
15239 => "000001",
15367 => "000001",
15495 => "000001",
15623 => "000001",
15751 => "000001",
15879 => "000001",
16007 => "000001",
16135 => "000001",
16263 => "000001",
13 => "000001",
141 => "000001",
269 => "000001",
397 => "000001",
525 => "000001",
653 => "000001",
781 => "000001",
909 => "000001",
1037 => "000001",
1165 => "000001",
1293 => "000001",
1421 => "000001",
1549 => "000001",
1677 => "000001",
1805 => "000001",
1933 => "000001",
2061 => "000001",
2189 => "000001",
2317 => "000001",
2445 => "000001",
2573 => "000001",
2701 => "000001",
2829 => "000001",
2957 => "000001",
3085 => "000001",
3213 => "000001",
3341 => "000001",
3469 => "000001",
3597 => "000001",
3725 => "000001",
3853 => "000001",
3981 => "000001",
4109 => "000001",
4237 => "000001",
4365 => "000001",
4493 => "000001",
4621 => "000001",
4749 => "000001",
4877 => "000001",
5005 => "000001",
5133 => "000001",
5261 => "000001",
5389 => "000001",
5517 => "000001",
5645 => "000001",
5773 => "000001",
5901 => "000001",
6029 => "000001",
6157 => "000001",
6285 => "000001",
6413 => "000001",
6541 => "000001",
6669 => "000001",
6797 => "000001",
6925 => "000001",
7053 => "000001",
7181 => "000001",
7309 => "000001",
7437 => "000001",
7565 => "000001",
7693 => "000001",
7821 => "000001",
7949 => "000001",
8077 => "000001",
8205 => "000001",
8333 => "000001",
8461 => "000001",
8589 => "000001",
8717 => "000001",
8845 => "000001",
8973 => "000001",
9101 => "000001",
9229 => "000001",
9357 => "000001",
9485 => "000001",
9613 => "000001",
9741 => "000001",
9869 => "000001",
9997 => "000001",
10125 => "000001",
10253 => "000001",
10381 => "000001",
10509 => "000001",
10637 => "000001",
10765 => "000001",
10893 => "000001",
11021 => "000001",
11149 => "000001",
11277 => "000001",
11405 => "000001",
11533 => "000001",
11661 => "000001",
11789 => "000001",
11917 => "000001",
12045 => "000001",
12173 => "000001",
12301 => "000001",
12429 => "000001",
12557 => "000001",
12685 => "000001",
12813 => "000001",
12941 => "000001",
13069 => "000001",
13197 => "000001",
13325 => "000001",
13453 => "000001",
13581 => "000001",
13709 => "000001",
13837 => "000001",
13965 => "000001",
14093 => "000001",
14221 => "000001",
14349 => "000001",
14477 => "000001",
14605 => "000001",
14733 => "000001",
14861 => "000001",
14989 => "000001",
15117 => "000001",
15245 => "000001",
15373 => "000001",
15501 => "000001",
15629 => "000001",
15757 => "000001",
15885 => "000001",
16013 => "000001",
16141 => "000001",
16269 => "000001",
19 => "000001",
147 => "000001",
275 => "000001",
403 => "000001",
531 => "000001",
659 => "000001",
787 => "000001",
915 => "000001",
1043 => "000001",
1171 => "000001",
1299 => "000001",
1427 => "000001",
1555 => "000001",
1683 => "000001",
1811 => "000001",
1939 => "000001",
2067 => "000001",
2195 => "000001",
2323 => "000001",
2451 => "000001",
2579 => "000001",
2707 => "000001",
2835 => "000001",
2963 => "000001",
3091 => "000001",
3219 => "000001",
3347 => "000001",
3475 => "000001",
3603 => "000001",
3731 => "000001",
3859 => "000001",
3987 => "000001",
4115 => "000001",
4243 => "000001",
4371 => "000001",
4499 => "000001",
4627 => "000001",
4755 => "000001",
4883 => "000001",
5011 => "000001",
5139 => "000001",
5267 => "000001",
5395 => "000001",
5523 => "000001",
5651 => "000001",
5779 => "000001",
5907 => "000001",
6035 => "000001",
6163 => "000001",
6291 => "000001",
6419 => "000001",
6547 => "000001",
6675 => "000001",
6803 => "000001",
6931 => "000001",
7059 => "000001",
7187 => "000001",
7315 => "000001",
7443 => "000001",
7571 => "000001",
7699 => "000001",
7827 => "000001",
7955 => "000001",
8083 => "000001",
8211 => "000001",
8339 => "000001",
8467 => "000001",
8595 => "000001",
8723 => "000001",
8851 => "000001",
8979 => "000001",
9107 => "000001",
9235 => "000001",
9363 => "000001",
9491 => "000001",
9619 => "000001",
9747 => "000001",
9875 => "000001",
10003 => "000001",
10131 => "000001",
10259 => "000001",
10387 => "000001",
10515 => "000001",
10643 => "000001",
10771 => "000001",
10899 => "000001",
11027 => "000001",
11155 => "000001",
11283 => "000001",
11411 => "000001",
11539 => "000001",
11667 => "000001",
11795 => "000001",
11923 => "000001",
12051 => "000001",
12179 => "000001",
12307 => "000001",
12435 => "000001",
12563 => "000001",
12691 => "000001",
12819 => "000001",
12947 => "000001",
13075 => "000001",
13203 => "000001",
13331 => "000001",
13459 => "000001",
13587 => "000001",
13715 => "000001",
13843 => "000001",
13971 => "000001",
14099 => "000001",
14227 => "000001",
14355 => "000001",
14483 => "000001",
14611 => "000001",
14739 => "000001",
14867 => "000001",
14995 => "000001",
15123 => "000001",
15251 => "000001",
15379 => "000001",
15507 => "000001",
15635 => "000001",
15763 => "000001",
15891 => "000001",
16019 => "000001",
16147 => "000001",
16275 => "000001",
25 => "000001",
153 => "000001",
281 => "000001",
409 => "000001",
537 => "000001",
665 => "000001",
793 => "000001",
921 => "000001",
1049 => "000001",
1177 => "000001",
1305 => "000001",
1433 => "000001",
1561 => "000001",
1689 => "000001",
1817 => "000001",
1945 => "000001",
2073 => "000001",
2201 => "000001",
2329 => "000001",
2457 => "000001",
2585 => "000001",
2713 => "000001",
2841 => "000001",
2969 => "000001",
3097 => "000001",
3225 => "000001",
3353 => "000001",
3481 => "000001",
3609 => "000001",
3737 => "000001",
3865 => "000001",
3993 => "000001",
4121 => "000001",
4249 => "000001",
4377 => "000001",
4505 => "000001",
4633 => "000001",
4761 => "000001",
4889 => "000001",
5017 => "000001",
5145 => "000001",
5273 => "000001",
5401 => "000001",
5529 => "000001",
5657 => "000001",
5785 => "000001",
5913 => "000001",
6041 => "000001",
6169 => "000001",
6297 => "000001",
6425 => "000001",
6553 => "000001",
6681 => "000001",
6809 => "000001",
6937 => "000001",
7065 => "000001",
7193 => "000001",
7321 => "000001",
7449 => "000001",
7577 => "000001",
7705 => "000001",
7833 => "000001",
7961 => "000001",
8089 => "000001",
8217 => "000001",
8345 => "000001",
8473 => "000001",
8601 => "000001",
8729 => "000001",
8857 => "000001",
8985 => "000001",
9113 => "000001",
9241 => "000001",
9369 => "000001",
9497 => "000001",
9625 => "000001",
9753 => "000001",
9881 => "000001",
10009 => "000001",
10137 => "000001",
10265 => "000001",
10393 => "000001",
10521 => "000001",
10649 => "000001",
10777 => "000001",
10905 => "000001",
11033 => "000001",
11161 => "000001",
11289 => "000001",
11417 => "000001",
11545 => "000001",
11673 => "000001",
11801 => "000001",
11929 => "000001",
12057 => "000001",
12185 => "000001",
12313 => "000001",
12441 => "000001",
12569 => "000001",
12697 => "000001",
12825 => "000001",
12953 => "000001",
13081 => "000001",
13209 => "000001",
13337 => "000001",
13465 => "000001",
13593 => "000001",
13721 => "000001",
13849 => "000001",
13977 => "000001",
14105 => "000001",
14233 => "000001",
14361 => "000001",
14489 => "000001",
14617 => "000001",
14745 => "000001",
14873 => "000001",
15001 => "000001",
15129 => "000001",
15257 => "000001",
15385 => "000001",
15513 => "000001",
15641 => "000001",
15769 => "000001",
15897 => "000001",
16025 => "000001",
16153 => "000001",
16281 => "000001",
31 => "000001",
159 => "000001",
287 => "000001",
415 => "000001",
543 => "000001",
671 => "000001",
799 => "000001",
927 => "000001",
1055 => "000001",
1183 => "000001",
1311 => "000001",
1439 => "000001",
1567 => "000001",
1695 => "000001",
1823 => "000001",
1951 => "000001",
2079 => "000001",
2207 => "000001",
2335 => "000001",
2463 => "000001",
2591 => "000001",
2719 => "000001",
2847 => "000001",
2975 => "000001",
3103 => "000001",
3231 => "000001",
3359 => "000001",
3487 => "000001",
3615 => "000001",
3743 => "000001",
3871 => "000001",
3999 => "000001",
4127 => "000001",
4255 => "000001",
4383 => "000001",
4511 => "000001",
4639 => "000001",
4767 => "000001",
4895 => "000001",
5023 => "000001",
5151 => "000001",
5279 => "000001",
5407 => "000001",
5535 => "000001",
5663 => "000001",
5791 => "000001",
5919 => "000001",
6047 => "000001",
6175 => "000001",
6303 => "000001",
6431 => "000001",
6559 => "000001",
6687 => "000001",
6815 => "000001",
6943 => "000001",
7071 => "000001",
7199 => "000001",
7327 => "000001",
7455 => "000001",
7583 => "000001",
7711 => "000001",
7839 => "000001",
7967 => "000001",
8095 => "000001",
8223 => "000001",
8351 => "000001",
8479 => "000001",
8607 => "000001",
8735 => "000001",
8863 => "000001",
8991 => "000001",
9119 => "000001",
9247 => "000001",
9375 => "000001",
9503 => "000001",
9631 => "000001",
9759 => "000001",
9887 => "000001",
10015 => "000001",
10143 => "000001",
10271 => "000001",
10399 => "000001",
10527 => "000001",
10655 => "000001",
10783 => "000001",
10911 => "000001",
11039 => "000001",
11167 => "000001",
11295 => "000001",
11423 => "000001",
11551 => "000001",
11679 => "000001",
11807 => "000001",
11935 => "000001",
12063 => "000001",
12191 => "000001",
12319 => "000001",
12447 => "000001",
12575 => "000001",
12703 => "000001",
12831 => "000001",
12959 => "000001",
13087 => "000001",
13215 => "000001",
13343 => "000001",
13471 => "000001",
13599 => "000001",
13727 => "000001",
13855 => "000001",
13983 => "000001",
14111 => "000001",
14239 => "000001",
14367 => "000001",
14495 => "000001",
14623 => "000001",
14751 => "000001",
14879 => "000001",
15007 => "000001",
15135 => "000001",
15263 => "000001",
15391 => "000001",
15519 => "000001",
15647 => "000001",
15775 => "000001",
15903 => "000001",
16031 => "000001",
16159 => "000001",
16287 => "000001",
37 => "000001",
165 => "000001",
293 => "000001",
421 => "000001",
549 => "000001",
677 => "000001",
805 => "000001",
933 => "000001",
1061 => "000001",
1189 => "000001",
1317 => "000001",
1445 => "000001",
1573 => "000001",
1701 => "000001",
1829 => "000001",
1957 => "000001",
2085 => "000001",
2213 => "000001",
2341 => "000001",
2469 => "000001",
2597 => "000001",
2725 => "000001",
2853 => "000001",
2981 => "000001",
3109 => "000001",
3237 => "000001",
3365 => "000001",
3493 => "000001",
3621 => "000001",
3749 => "000001",
3877 => "000001",
4005 => "000001",
4133 => "000001",
4261 => "000001",
4389 => "000001",
4517 => "000001",
4645 => "000001",
4773 => "000001",
4901 => "000001",
5029 => "000001",
5157 => "000001",
5285 => "000001",
5413 => "000001",
5541 => "000001",
5669 => "000001",
5797 => "000001",
5925 => "000001",
6053 => "000001",
6181 => "000001",
6309 => "000001",
6437 => "000001",
6565 => "000001",
6693 => "000001",
6821 => "000001",
6949 => "000001",
7077 => "000001",
7205 => "000001",
7333 => "000001",
7461 => "000001",
7589 => "000001",
7717 => "000001",
7845 => "000001",
7973 => "000001",
8101 => "000001",
8229 => "000001",
8357 => "000001",
8485 => "000001",
8613 => "000001",
8741 => "000001",
8869 => "000001",
8997 => "000001",
9125 => "000001",
9253 => "000001",
9381 => "000001",
9509 => "000001",
9637 => "000001",
9765 => "000001",
9893 => "000001",
10021 => "000001",
10149 => "000001",
10277 => "000001",
10405 => "000001",
10533 => "000001",
10661 => "000001",
10789 => "000001",
10917 => "000001",
11045 => "000001",
11173 => "000001",
11301 => "000001",
11429 => "000001",
11557 => "000001",
11685 => "000001",
11813 => "000001",
11941 => "000001",
12069 => "000001",
12197 => "000001",
12325 => "000001",
12453 => "000001",
12581 => "000001",
12709 => "000001",
12837 => "000001",
12965 => "000001",
13093 => "000001",
13221 => "000001",
13349 => "000001",
13477 => "000001",
13605 => "000001",
13733 => "000001",
13861 => "000001",
13989 => "000001",
14117 => "000001",
14245 => "000001",
14373 => "000001",
14501 => "000001",
14629 => "000001",
14757 => "000001",
14885 => "000001",
15013 => "000001",
15141 => "000001",
15269 => "000001",
15397 => "000001",
15525 => "000001",
15653 => "000001",
15781 => "000001",
15909 => "000001",
16037 => "000001",
16165 => "000001",
16293 => "000001",
43 => "000001",
171 => "000001",
299 => "000001",
427 => "000001",
555 => "000001",
683 => "000001",
811 => "000001",
939 => "000001",
1067 => "000001",
1195 => "000001",
1323 => "000001",
1451 => "000001",
1579 => "000001",
1707 => "000001",
1835 => "000001",
1963 => "000001",
2091 => "000001",
2219 => "000001",
2347 => "000001",
2475 => "000001",
2603 => "000001",
2731 => "000001",
2859 => "000001",
2987 => "000001",
3115 => "000001",
3243 => "000001",
3371 => "000001",
3499 => "000001",
3627 => "000001",
3755 => "000001",
3883 => "000001",
4011 => "000001",
4139 => "000001",
4267 => "000001",
4395 => "000001",
4523 => "000001",
4651 => "000001",
4779 => "000001",
4907 => "000001",
5035 => "000001",
5163 => "000001",
5291 => "000001",
5419 => "000001",
5547 => "000001",
5675 => "000001",
5803 => "000001",
5931 => "000001",
6059 => "000001",
6187 => "000001",
6315 => "000001",
6443 => "000001",
6571 => "000001",
6699 => "000001",
6827 => "000001",
6955 => "000001",
7083 => "000001",
7211 => "000001",
7339 => "000001",
7467 => "000001",
7595 => "000001",
7723 => "000001",
7851 => "000001",
7979 => "000001",
8107 => "000001",
8235 => "000001",
8363 => "000001",
8491 => "000001",
8619 => "000001",
8747 => "000001",
8875 => "000001",
9003 => "000001",
9131 => "000001",
9259 => "000001",
9387 => "000001",
9515 => "000001",
9643 => "000001",
9771 => "000001",
9899 => "000001",
10027 => "000001",
10155 => "000001",
10283 => "000001",
10411 => "000001",
10539 => "000001",
10667 => "000001",
10795 => "000001",
10923 => "000001",
11051 => "000001",
11179 => "000001",
11307 => "000001",
11435 => "000001",
11563 => "000001",
11691 => "000001",
11819 => "000001",
11947 => "000001",
12075 => "000001",
12203 => "000001",
12331 => "000001",
12459 => "000001",
12587 => "000001",
12715 => "000001",
12843 => "000001",
12971 => "000001",
13099 => "000001",
13227 => "000001",
13355 => "000001",
13483 => "000001",
13611 => "000001",
13739 => "000001",
13867 => "000001",
13995 => "000001",
14123 => "000001",
14251 => "000001",
14379 => "000001",
14507 => "000001",
14635 => "000001",
14763 => "000001",
14891 => "000001",
15019 => "000001",
15147 => "000001",
15275 => "000001",
15403 => "000001",
15531 => "000001",
15659 => "000001",
15787 => "000001",
15915 => "000001",
16043 => "000001",
16171 => "000001",
16299 => "000001",
49 => "000001",
177 => "000001",
305 => "000001",
433 => "000001",
561 => "000001",
689 => "000001",
817 => "000001",
945 => "000001",
1073 => "000001",
1201 => "000001",
1329 => "000001",
1457 => "000001",
1585 => "000001",
1713 => "000001",
1841 => "000001",
1969 => "000001",
2097 => "000001",
2225 => "000001",
2353 => "000001",
2481 => "000001",
2609 => "000001",
2737 => "000001",
2865 => "000001",
2993 => "000001",
3121 => "000001",
3249 => "000001",
3377 => "000001",
3505 => "000001",
3633 => "000001",
3761 => "000001",
3889 => "000001",
4017 => "000001",
4145 => "000001",
4273 => "000001",
4401 => "000001",
4529 => "000001",
4657 => "000001",
4785 => "000001",
4913 => "000001",
5041 => "000001",
5169 => "000001",
5297 => "000001",
5425 => "000001",
5553 => "000001",
5681 => "000001",
5809 => "000001",
5937 => "000001",
6065 => "000001",
6193 => "000001",
6321 => "000001",
6449 => "000001",
6577 => "000001",
6705 => "000001",
6833 => "000001",
6961 => "000001",
7089 => "000001",
7217 => "000001",
7345 => "000001",
7473 => "000001",
7601 => "000001",
7729 => "000001",
7857 => "000001",
7985 => "000001",
8113 => "000001",
8241 => "000001",
8369 => "000001",
8497 => "000001",
8625 => "000001",
8753 => "000001",
8881 => "000001",
9009 => "000001",
9137 => "000001",
9265 => "000001",
9393 => "000001",
9521 => "000001",
9649 => "000001",
9777 => "000001",
9905 => "000001",
10033 => "000001",
10161 => "000001",
10289 => "000001",
10417 => "000001",
10545 => "000001",
10673 => "000001",
10801 => "000001",
10929 => "000001",
11057 => "000001",
11185 => "000001",
11313 => "000001",
11441 => "000001",
11569 => "000001",
11697 => "000001",
11825 => "000001",
11953 => "000001",
12081 => "000001",
12209 => "000001",
12337 => "000001",
12465 => "000001",
12593 => "000001",
12721 => "000001",
12849 => "000001",
12977 => "000001",
13105 => "000001",
13233 => "000001",
13361 => "000001",
13489 => "000001",
13617 => "000001",
13745 => "000001",
13873 => "000001",
14001 => "000001",
14129 => "000001",
14257 => "000001",
14385 => "000001",
14513 => "000001",
14641 => "000001",
14769 => "000001",
14897 => "000001",
15025 => "000001",
15153 => "000001",
15281 => "000001",
15409 => "000001",
15537 => "000001",
15665 => "000001",
15793 => "000001",
15921 => "000001",
16049 => "000001",
16177 => "000001",
16305 => "000001",
55 => "000001",
183 => "000001",
311 => "000001",
439 => "000001",
567 => "000001",
695 => "000001",
823 => "000001",
951 => "000001",
1079 => "000001",
1207 => "000001",
1335 => "000001",
1463 => "000001",
1591 => "000001",
1719 => "000001",
1847 => "000001",
1975 => "000001",
2103 => "000001",
2231 => "000001",
2359 => "000001",
2487 => "000001",
2615 => "000001",
2743 => "000001",
2871 => "000001",
2999 => "000001",
3127 => "000001",
3255 => "000001",
3383 => "000001",
3511 => "000001",
3639 => "000001",
3767 => "000001",
3895 => "000001",
4023 => "000001",
4151 => "000001",
4279 => "000001",
4407 => "000001",
4535 => "000001",
4663 => "000001",
4791 => "000001",
4919 => "000001",
5047 => "000001",
5175 => "000001",
5303 => "000001",
5431 => "000001",
5559 => "000001",
5687 => "000001",
5815 => "000001",
5943 => "000001",
6071 => "000001",
6199 => "000001",
6327 => "000001",
6455 => "000001",
6583 => "000001",
6711 => "000001",
6839 => "000001",
6967 => "000001",
7095 => "000001",
7223 => "000001",
7351 => "000001",
7479 => "000001",
7607 => "000001",
7735 => "000001",
7863 => "000001",
7991 => "000001",
8119 => "000001",
8247 => "000001",
8375 => "000001",
8503 => "000001",
8631 => "000001",
8759 => "000001",
8887 => "000001",
9015 => "000001",
9143 => "000001",
9271 => "000001",
9399 => "000001",
9527 => "000001",
9655 => "000001",
9783 => "000001",
9911 => "000001",
10039 => "000001",
10167 => "000001",
10295 => "000001",
10423 => "000001",
10551 => "000001",
10679 => "000001",
10807 => "000001",
10935 => "000001",
11063 => "000001",
11191 => "000001",
11319 => "000001",
11447 => "000001",
11575 => "000001",
11703 => "000001",
11831 => "000001",
11959 => "000001",
12087 => "000001",
12215 => "000001",
12343 => "000001",
12471 => "000001",
12599 => "000001",
12727 => "000001",
12855 => "000001",
12983 => "000001",
13111 => "000001",
13239 => "000001",
13367 => "000001",
13495 => "000001",
13623 => "000001",
13751 => "000001",
13879 => "000001",
14007 => "000001",
14135 => "000001",
14263 => "000001",
14391 => "000001",
14519 => "000001",
14647 => "000001",
14775 => "000001",
14903 => "000001",
15031 => "000001",
15159 => "000001",
15287 => "000001",
15415 => "000001",
15543 => "000001",
15671 => "000001",
15799 => "000001",
15927 => "000001",
16055 => "000001",
16183 => "000001",
16311 => "000001",
61 => "000001",
189 => "000001",
317 => "000001",
445 => "000001",
573 => "000001",
701 => "000001",
829 => "000001",
957 => "000001",
1085 => "000001",
1213 => "000001",
1341 => "000001",
1469 => "000001",
1597 => "000001",
1725 => "000001",
1853 => "000001",
1981 => "000001",
2109 => "000001",
2237 => "000001",
2365 => "000001",
2493 => "000001",
2621 => "000001",
2749 => "000001",
2877 => "000001",
3005 => "000001",
3133 => "000001",
3261 => "000001",
3389 => "000001",
3517 => "000001",
3645 => "000001",
3773 => "000001",
3901 => "000001",
4029 => "000001",
4157 => "000001",
4285 => "000001",
4413 => "000001",
4541 => "000001",
4669 => "000001",
4797 => "000001",
4925 => "000001",
5053 => "000001",
5181 => "000001",
5309 => "000001",
5437 => "000001",
5565 => "000001",
5693 => "000001",
5821 => "000001",
5949 => "000001",
6077 => "000001",
6205 => "000001",
6333 => "000001",
6461 => "000001",
6589 => "000001",
6717 => "000001",
6845 => "000001",
6973 => "000001",
7101 => "000001",
7229 => "000001",
7357 => "000001",
7485 => "000001",
7613 => "000001",
7741 => "000001",
7869 => "000001",
7997 => "000001",
8125 => "000001",
8253 => "000001",
8381 => "000001",
8509 => "000001",
8637 => "000001",
8765 => "000001",
8893 => "000001",
9021 => "000001",
9149 => "000001",
9277 => "000001",
9405 => "000001",
9533 => "000001",
9661 => "000001",
9789 => "000001",
9917 => "000001",
10045 => "000001",
10173 => "000001",
10301 => "000001",
10429 => "000001",
10557 => "000001",
10685 => "000001",
10813 => "000001",
10941 => "000001",
11069 => "000001",
11197 => "000001",
11325 => "000001",
11453 => "000001",
11581 => "000001",
11709 => "000001",
11837 => "000001",
11965 => "000001",
12093 => "000001",
12221 => "000001",
12349 => "000001",
12477 => "000001",
12605 => "000001",
12733 => "000001",
12861 => "000001",
12989 => "000001",
13117 => "000001",
13245 => "000001",
13373 => "000001",
13501 => "000001",
13629 => "000001",
13757 => "000001",
13885 => "000001",
14013 => "000001",
14141 => "000001",
14269 => "000001",
14397 => "000001",
14525 => "000001",
14653 => "000001",
14781 => "000001",
14909 => "000001",
15037 => "000001",
15165 => "000001",
15293 => "000001",
15421 => "000001",
15549 => "000001",
15677 => "000001",
15805 => "000001",
15933 => "000001",
16061 => "000001",
16189 => "000001",
16317 => "000001",
67 => "000001",
195 => "000001",
323 => "000001",
451 => "000001",
579 => "000001",
707 => "000001",
835 => "000001",
963 => "000001",
1091 => "000001",
1219 => "000001",
1347 => "000001",
1475 => "000001",
1603 => "000001",
1731 => "000001",
1859 => "000001",
1987 => "000001",
2115 => "000001",
2243 => "000001",
2371 => "000001",
2499 => "000001",
2627 => "000001",
2755 => "000001",
2883 => "000001",
3011 => "000001",
3139 => "000001",
3267 => "000001",
3395 => "000001",
3523 => "000001",
3651 => "000001",
3779 => "000001",
3907 => "000001",
4035 => "000001",
4163 => "000001",
4291 => "000001",
4419 => "000001",
4547 => "000001",
4675 => "000001",
4803 => "000001",
4931 => "000001",
5059 => "000001",
5187 => "000001",
5315 => "000001",
5443 => "000001",
5571 => "000001",
5699 => "000001",
5827 => "000001",
5955 => "000001",
6083 => "000001",
6211 => "000001",
6339 => "000001",
6467 => "000001",
6595 => "000001",
6723 => "000001",
6851 => "000001",
6979 => "000001",
7107 => "000001",
7235 => "000001",
7363 => "000001",
7491 => "000001",
7619 => "000001",
7747 => "000001",
7875 => "000001",
8003 => "000001",
8131 => "000001",
8259 => "000001",
8387 => "000001",
8515 => "000001",
8643 => "000001",
8771 => "000001",
8899 => "000001",
9027 => "000001",
9155 => "000001",
9283 => "000001",
9411 => "000001",
9539 => "000001",
9667 => "000001",
9795 => "000001",
9923 => "000001",
10051 => "000001",
10179 => "000001",
10307 => "000001",
10435 => "000001",
10563 => "000001",
10691 => "000001",
10819 => "000001",
10947 => "000001",
11075 => "000001",
11203 => "000001",
11331 => "000001",
11459 => "000001",
11587 => "000001",
11715 => "000001",
11843 => "000001",
11971 => "000001",
12099 => "000001",
12227 => "000001",
12355 => "000001",
12483 => "000001",
12611 => "000001",
12739 => "000001",
12867 => "000001",
12995 => "000001",
13123 => "000001",
13251 => "000001",
13379 => "000001",
13507 => "000001",
13635 => "000001",
13763 => "000001",
13891 => "000001",
14019 => "000001",
14147 => "000001",
14275 => "000001",
14403 => "000001",
14531 => "000001",
14659 => "000001",
14787 => "000001",
14915 => "000001",
15043 => "000001",
15171 => "000001",
15299 => "000001",
15427 => "000001",
15555 => "000001",
15683 => "000001",
15811 => "000001",
15939 => "000001",
16067 => "000001",
16195 => "000001",
16323 => "000001",
73 => "000001",
201 => "000001",
329 => "000001",
457 => "000001",
585 => "000001",
713 => "000001",
841 => "000001",
969 => "000001",
1097 => "000001",
1225 => "000001",
1353 => "000001",
1481 => "000001",
1609 => "000001",
1737 => "000001",
1865 => "000001",
1993 => "000001",
2121 => "000001",
2249 => "000001",
2377 => "000001",
2505 => "000001",
2633 => "000001",
2761 => "000001",
2889 => "000001",
3017 => "000001",
3145 => "000001",
3273 => "000001",
3401 => "000001",
3529 => "000001",
3657 => "000001",
3785 => "000001",
3913 => "000001",
4041 => "000001",
4169 => "000001",
4297 => "000001",
4425 => "000001",
4553 => "000001",
4681 => "000001",
4809 => "000001",
4937 => "000001",
5065 => "000001",
5193 => "000001",
5321 => "000001",
5449 => "000001",
5577 => "000001",
5705 => "000001",
5833 => "000001",
5961 => "000001",
6089 => "000001",
6217 => "000001",
6345 => "000001",
6473 => "000001",
6601 => "000001",
6729 => "000001",
6857 => "000001",
6985 => "000001",
7113 => "000001",
7241 => "000001",
7369 => "000001",
7497 => "000001",
7625 => "000001",
7753 => "000001",
7881 => "000001",
8009 => "000001",
8137 => "000001",
8265 => "000001",
8393 => "000001",
8521 => "000001",
8649 => "000001",
8777 => "000001",
8905 => "000001",
9033 => "000001",
9161 => "000001",
9289 => "000001",
9417 => "000001",
9545 => "000001",
9673 => "000001",
9801 => "000001",
9929 => "000001",
10057 => "000001",
10185 => "000001",
10313 => "000001",
10441 => "000001",
10569 => "000001",
10697 => "000001",
10825 => "000001",
10953 => "000001",
11081 => "000001",
11209 => "000001",
11337 => "000001",
11465 => "000001",
11593 => "000001",
11721 => "000001",
11849 => "000001",
11977 => "000001",
12105 => "000001",
12233 => "000001",
12361 => "000001",
12489 => "000001",
12617 => "000001",
12745 => "000001",
12873 => "000001",
13001 => "000001",
13129 => "000001",
13257 => "000001",
13385 => "000001",
13513 => "000001",
13641 => "000001",
13769 => "000001",
13897 => "000001",
14025 => "000001",
14153 => "000001",
14281 => "000001",
14409 => "000001",
14537 => "000001",
14665 => "000001",
14793 => "000001",
14921 => "000001",
15049 => "000001",
15177 => "000001",
15305 => "000001",
15433 => "000001",
15561 => "000001",
15689 => "000001",
15817 => "000001",
15945 => "000001",
16073 => "000001",
16201 => "000001",
16329 => "000001",
79 => "000010",
207 => "000010",
335 => "000010",
463 => "000010",
591 => "000010",
719 => "000010",
847 => "000010",
975 => "000010",
1103 => "000010",
1231 => "000010",
1359 => "000010",
1487 => "000010",
1615 => "000010",
1743 => "000010",
1871 => "000010",
1999 => "000010",
2127 => "000010",
2255 => "000010",
2383 => "000010",
2511 => "000010",
2639 => "000010",
2767 => "000010",
2895 => "000010",
3023 => "000010",
3151 => "000010",
3279 => "000010",
3407 => "000010",
3535 => "000010",
3663 => "000010",
3791 => "000010",
3919 => "000010",
4047 => "000010",
4175 => "000010",
4303 => "000010",
4431 => "000010",
4559 => "000010",
4687 => "000010",
4815 => "000010",
4943 => "000010",
5071 => "000010",
5199 => "000010",
5327 => "000010",
5455 => "000010",
5583 => "000010",
5711 => "000010",
5839 => "000010",
5967 => "000010",
6095 => "000010",
6223 => "000010",
6351 => "000010",
6479 => "000010",
6607 => "000010",
6735 => "000010",
6863 => "000010",
6991 => "000010",
7119 => "000010",
7247 => "000010",
7375 => "000010",
7503 => "000010",
7631 => "000010",
7759 => "000010",
7887 => "000010",
8015 => "000010",
8143 => "000010",
8271 => "000010",
8399 => "000010",
8527 => "000010",
8655 => "000010",
8783 => "000010",
8911 => "000010",
9039 => "000010",
9167 => "000010",
9295 => "000010",
9423 => "000010",
9551 => "000010",
9679 => "000010",
9807 => "000010",
9935 => "000010",
10063 => "000010",
10191 => "000010",
10319 => "000010",
10447 => "000010",
10575 => "000010",
10703 => "000010",
10831 => "000010",
10959 => "000010",
11087 => "000010",
11215 => "000010",
11343 => "000010",
11471 => "000010",
11599 => "000010",
11727 => "000010",
11855 => "000010",
11983 => "000010",
12111 => "000010",
12239 => "000010",
12367 => "000010",
12495 => "000010",
12623 => "000010",
12751 => "000010",
12879 => "000010",
13007 => "000010",
13135 => "000010",
13263 => "000010",
13391 => "000010",
13519 => "000010",
13647 => "000010",
13775 => "000010",
13903 => "000010",
14031 => "000010",
14159 => "000010",
14287 => "000010",
14415 => "000010",
14543 => "000010",
14671 => "000010",
14799 => "000010",
14927 => "000010",
15055 => "000010",
15183 => "000010",
15311 => "000010",
15439 => "000010",
15567 => "000010",
15695 => "000010",
15823 => "000010",
15951 => "000010",
16079 => "000010",
16207 => "000010",
16335 => "000010",


    others => (others => '0')
    );

    attribute ram_style : string;
    attribute ram_style of tile_data_map : signal is "block";
    

begin

    -- Compute tile index from view position
    s_view_index(13 downto 7) <= i_view_y(9 downto 3);
    s_view_index(6 downto 0)  <= i_view_x(9 downto 3);

    -- Read output values
    o_tile_id <= tile_data_map(to_integer(unsigned(s_view_index)))(4 downto 0);
    o_flip_y  <= tile_data_map(to_integer(unsigned(s_view_index)))(5);
    o_pix_x   <= i_view_x(2 downto 0);
    o_pix_y   <= i_view_y(2 downto 0);

    -- Write process
    process(i_clk)
        variable write_index : std_logic_vector(13 downto 0);
        variable new_data    : std_logic_vector(5 downto 0);
    begin
        if rising_edge(i_clk) then
            if (i_ch_we_tileBack = '1') then
                write_index := i_row & i_col;
                new_data := tile_data_map(to_integer(unsigned(write_index)));

                -- Update tile_id if required
                if i_ch_tile_id = '1' then
                    new_data(4 downto 0) := i_tile_id;
                end if;

                -- Update flip_y if required
                if i_ch_flipY = '1' then
                    new_data(5) := i_flip_y;
                end if;

                -- Write back to BRAM
                tile_data_map(to_integer(unsigned(write_index))) <= new_data;
            end if;
        end if;
    end process;

end Behavioral;
