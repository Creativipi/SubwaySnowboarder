----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08.06.2025 00:00:57
-- Design Name: 
-- Module Name: ActorMgmt - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
 
 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
 
-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
 
entity ActorMgmt is
    Port (
        -- Position du pixel dans le viewport
        i_view_x : in STD_LOGIC_VECTOR (9 downto 0);
        i_view_y : in STD_LOGIC_VECTOR (9 downto 0);
 
        -- Mise ? jour des acteurs (position RELATIVE AU VIEWPORT)
        i_act_id : in STD_LOGIC_VECTOR (2 downto 0);
        i_newpos_x : in STD_LOGIC_VECTOR (9 downto 0);
        i_newpos_y : in STD_LOGIC_VECTOR (9 downto 0);
        i_tile_id : in STD_LOGIC_VECTOR (3 downto 0);
        i_flip_x : in STD_LOGIC;
        i_flip_y : in STD_LOGIC;
        i_ch_setpos : in STD_LOGIC;
        i_ch_tile_id : in STD_LOGIC;
        i_ch_flipX : in STD_LOGIC;
        i_ch_flipY : in STD_LOGIC;
        i_clk : in STD_LOGIC;
        i_ch_x : in std_logic_vector (3 downto 0);
        i_ch_y : in std_logic_vector (3 downto 0);
        i_ch_cc : in std_logic_vector (3 downto 0);
        i_tile_id_write : in std_logic_vector (3 downto 0);
        i_ch_we : in std_logic;
 
        -- R?sultat : info du pixel
        o_tile_id : out STD_LOGIC_VECTOR (3 downto 0);
        o_flip_x : out STD_LOGIC;
        o_flip_y : out STD_LOGIC;
        o_pix_x : out STD_LOGIC_VECTOR (3 downto 0);
        o_pix_y : out STD_LOGIC_VECTOR (3 downto 0);
        o_is_actor_present : out STD_LOGIC
    );
end ActorMgmt;
 
architecture Behavioral of ActorMgmt is
    -- Sparse array de 8 acteurs
    type pos_array_t is array (0 to 7) of std_logic_vector(9 downto 0);
    type tile_array_t is array (0 to 7) of std_logic_vector(3 downto 0);
    type flip_array_t is array (0 to 7) of std_logic;
 
    signal actor_pos_x : pos_array_t := (
    0 => std_logic_vector(to_unsigned(320, 10)), -- acteur 0 au centre du viewport
    1 => std_logic_vector(to_unsigned(336, 10)), -- acteur 1 juste ? droite (16 px)
    others => (others => '0')
);
 
signal actor_pos_y : pos_array_t := (
    0 => std_logic_vector(to_unsigned(180, 10)), -- centr? verticalement
    1 => std_logic_vector(to_unsigned(180, 10)),
    others => (others => '0')
);
 
signal actor_tile_id : tile_array_t := (
    others => std_logic_vector(to_unsigned(0, 4))
);
 
    signal actor_flip_x : flip_array_t := (others => '0');
    signal actor_flip_y : flip_array_t := (others => '0');
 
    signal s_actor_hit : std_logic_vector(7 downto 0);
    signal s_found : std_logic;
    type tile_d_array_a is array (0 to 4095) of std_logic;
    signal tile_data_map_a : tile_d_array_a := (
    0 => '1',
1 => '1',
2 => '1',
3 => '1',
4 => '1',
5 => '1',
6 => '1',
7 => '1',
8 => '0',
9 => '1',
10 => '1',
11 => '1',
12 => '1',
13 => '1',
14 => '1',
15 => '1',
16 => '1',
17 => '1',
18 => '1',
19 => '1',
20 => '1',
21 => '1',
22 => '1',
23 => '0',
24 => '0',
25 => '1',
26 => '1',
27 => '1',
28 => '1',
29 => '1',
30 => '1',
31 => '1',
32 => '1',
33 => '1',
34 => '0',
35 => '1',
36 => '1',
37 => '1',
38 => '0',
39 => '0',
40 => '0',
41 => '1',
42 => '1',
43 => '1',
44 => '1',
45 => '1',
46 => '1',
47 => '1',
48 => '1',
49 => '0',
50 => '0',
51 => '0',
52 => '1',
53 => '0',
54 => '0',
55 => '0',
56 => '0',
57 => '1',
58 => '1',
59 => '1',
60 => '1',
61 => '1',
62 => '1',
63 => '1',
64 => '1',
65 => '0',
66 => '0',
67 => '0',
68 => '0',
69 => '0',
70 => '0',
71 => '0',
72 => '0',
73 => '1',
74 => '1',
75 => '1',
76 => '1',
77 => '1',
78 => '1',
79 => '1',
80 => '1',
81 => '1',
82 => '0',
83 => '0',
84 => '0',
85 => '0',
86 => '0',
87 => '0',
88 => '0',
89 => '1',
90 => '1',
91 => '1',
92 => '1',
93 => '1',
94 => '1',
95 => '1',
96 => '1',
97 => '1',
98 => '0',
99 => '0',
100 => '0',
101 => '0',
102 => '0',
103 => '0',
104 => '0',
105 => '1',
106 => '1',
107 => '1',
108 => '1',
109 => '1',
110 => '1',
111 => '1',
112 => '1',
113 => '0',
114 => '0',
115 => '0',
116 => '0',
117 => '0',
118 => '0',
119 => '0',
120 => '0',
121 => '0',
122 => '0',
123 => '0',
124 => '0',
125 => '0',
126 => '1',
127 => '0',
128 => '1',
129 => '0',
130 => '0',
131 => '0',
132 => '0',
133 => '0',
134 => '0',
135 => '0',
136 => '0',
137 => '0',
138 => '0',
139 => '0',
140 => '0',
141 => '0',
142 => '0',
143 => '1',
144 => '0',
145 => '0',
146 => '0',
147 => '0',
148 => '0',
149 => '0',
150 => '0',
151 => '0',
152 => '0',
153 => '0',
154 => '0',
155 => '0',
156 => '0',
157 => '0',
158 => '1',
159 => '1',
160 => '0',
161 => '0',
162 => '0',
163 => '0',
164 => '0',
165 => '0',
166 => '0',
167 => '0',
168 => '0',
169 => '0',
170 => '0',
171 => '0',
172 => '0',
173 => '1',
174 => '1',
175 => '1',
176 => '0',
177 => '0',
178 => '0',
179 => '0',
180 => '0',
181 => '0',
182 => '0',
183 => '0',
184 => '0',
185 => '0',
186 => '0',
187 => '0',
188 => '1',
189 => '1',
190 => '1',
191 => '1',
192 => '0',
193 => '0',
194 => '0',
195 => '0',
196 => '0',
197 => '0',
198 => '0',
199 => '0',
200 => '0',
201 => '0',
202 => '0',
203 => '1',
204 => '1',
205 => '1',
206 => '1',
207 => '1',
208 => '1',
209 => '0',
210 => '0',
211 => '0',
212 => '0',
213 => '0',
214 => '0',
215 => '0',
216 => '0',
217 => '0',
218 => '1',
219 => '1',
220 => '1',
221 => '1',
222 => '1',
223 => '1',
224 => '1',
225 => '1',
226 => '0',
227 => '0',
228 => '0',
229 => '0',
230 => '0',
231 => '0',
232 => '0',
233 => '1',
234 => '1',
235 => '1',
236 => '1',
237 => '1',
238 => '1',
239 => '1',
240 => '1',
241 => '1',
242 => '1',
243 => '0',
244 => '0',
245 => '0',
246 => '0',
247 => '1',
248 => '1',
249 => '1',
250 => '1',
251 => '1',
252 => '1',
253 => '1',
254 => '1',
255 => '1',
256 => '1',
257 => '1',
258 => '1',
259 => '1',
260 => '1',
261 => '1',
262 => '1',
263 => '1',
264 => '1',
265 => '0',
266 => '0',
267 => '0',
268 => '0',
269 => '1',
270 => '1',
271 => '0',
272 => '1',
273 => '1',
274 => '1',
275 => '1',
276 => '1',
277 => '1',
278 => '1',
279 => '0',
280 => '0',
281 => '0',
282 => '0',
283 => '0',
284 => '0',
285 => '0',
286 => '0',
287 => '0',
288 => '1',
289 => '1',
290 => '1',
291 => '1',
292 => '1',
293 => '1',
294 => '0',
295 => '0',
296 => '0',
297 => '0',
298 => '0',
299 => '0',
300 => '0',
301 => '0',
302 => '0',
303 => '0',
304 => '1',
305 => '1',
306 => '1',
307 => '1',
308 => '1',
309 => '0',
310 => '0',
311 => '0',
312 => '0',
313 => '0',
314 => '0',
315 => '0',
316 => '0',
317 => '0',
318 => '0',
319 => '0',
320 => '1',
321 => '1',
322 => '1',
323 => '1',
324 => '0',
325 => '0',
326 => '0',
327 => '0',
328 => '0',
329 => '0',
330 => '0',
331 => '0',
332 => '0',
333 => '0',
334 => '0',
335 => '0',
336 => '1',
337 => '1',
338 => '1',
339 => '0',
340 => '0',
341 => '0',
342 => '0',
343 => '0',
344 => '0',
345 => '0',
346 => '0',
347 => '0',
348 => '0',
349 => '0',
350 => '0',
351 => '0',
352 => '1',
353 => '1',
354 => '0',
355 => '0',
356 => '0',
357 => '0',
358 => '0',
359 => '0',
360 => '0',
361 => '0',
362 => '0',
363 => '0',
364 => '0',
365 => '0',
366 => '0',
367 => '0',
368 => '1',
369 => '0',
370 => '0',
371 => '0',
372 => '0',
373 => '0',
374 => '0',
375 => '0',
376 => '0',
377 => '0',
378 => '0',
379 => '0',
380 => '0',
381 => '0',
382 => '0',
383 => '0',
384 => '0',
385 => '0',
386 => '0',
387 => '0',
388 => '0',
389 => '0',
390 => '0',
391 => '0',
392 => '0',
393 => '0',
394 => '0',
395 => '0',
396 => '0',
397 => '0',
398 => '0',
399 => '1',
400 => '0',
401 => '0',
402 => '0',
403 => '0',
404 => '0',
405 => '0',
406 => '0',
407 => '0',
408 => '0',
409 => '0',
410 => '0',
411 => '0',
412 => '0',
413 => '0',
414 => '1',
415 => '1',
416 => '0',
417 => '0',
418 => '0',
419 => '0',
420 => '0',
421 => '0',
422 => '0',
423 => '0',
424 => '0',
425 => '0',
426 => '0',
427 => '0',
428 => '0',
429 => '1',
430 => '1',
431 => '1',
432 => '0',
433 => '0',
434 => '0',
435 => '0',
436 => '0',
437 => '0',
438 => '0',
439 => '0',
440 => '0',
441 => '0',
442 => '0',
443 => '0',
444 => '1',
445 => '1',
446 => '1',
447 => '1',
448 => '0',
449 => '0',
450 => '0',
451 => '0',
452 => '0',
453 => '0',
454 => '0',
455 => '0',
456 => '0',
457 => '0',
458 => '0',
459 => '1',
460 => '1',
461 => '1',
462 => '1',
463 => '1',
464 => '0',
465 => '0',
466 => '0',
467 => '0',
468 => '0',
469 => '0',
470 => '0',
471 => '0',
472 => '0',
473 => '0',
474 => '1',
475 => '1',
476 => '1',
477 => '1',
478 => '1',
479 => '1',
480 => '0',
481 => '0',
482 => '0',
483 => '0',
484 => '0',
485 => '0',
486 => '0',
487 => '0',
488 => '0',
489 => '1',
490 => '1',
491 => '1',
492 => '1',
493 => '1',
494 => '1',
495 => '1',
496 => '0',
497 => '0',
498 => '0',
499 => '0',
500 => '0',
501 => '0',
502 => '0',
503 => '0',
504 => '1',
505 => '1',
506 => '1',
507 => '1',
508 => '1',
509 => '1',
510 => '1',
511 => '1',
512 => '1',
513 => '1',
514 => '1',
515 => '1',
516 => '1',
517 => '1',
518 => '1',
519 => '0',
520 => '0',
521 => '1',
522 => '1',
523 => '1',
524 => '1',
525 => '1',
526 => '1',
527 => '1',
528 => '1',
529 => '1',
530 => '1',
531 => '1',
532 => '1',
533 => '1',
534 => '1',
535 => '0',
536 => '0',
537 => '0',
538 => '1',
539 => '1',
540 => '1',
541 => '1',
542 => '1',
543 => '1',
544 => '1',
545 => '1',
546 => '1',
547 => '1',
548 => '1',
549 => '1',
550 => '0',
551 => '0',
552 => '0',
553 => '0',
554 => '0',
555 => '1',
556 => '1',
557 => '1',
558 => '1',
559 => '1',
560 => '1',
561 => '1',
562 => '1',
563 => '1',
564 => '1',
565 => '0',
566 => '0',
567 => '0',
568 => '0',
569 => '0',
570 => '0',
571 => '0',
572 => '1',
573 => '1',
574 => '1',
575 => '1',
576 => '1',
577 => '1',
578 => '1',
579 => '1',
580 => '0',
581 => '0',
582 => '0',
583 => '0',
584 => '0',
585 => '0',
586 => '0',
587 => '0',
588 => '0',
589 => '1',
590 => '1',
591 => '1',
592 => '1',
593 => '1',
594 => '1',
595 => '1',
596 => '0',
597 => '0',
598 => '0',
599 => '0',
600 => '0',
601 => '0',
602 => '0',
603 => '0',
604 => '0',
605 => '1',
606 => '1',
607 => '1',
608 => '1',
609 => '1',
610 => '1',
611 => '0',
612 => '0',
613 => '0',
614 => '0',
615 => '0',
616 => '0',
617 => '0',
618 => '0',
619 => '0',
620 => '0',
621 => '0',
622 => '1',
623 => '1',
624 => '1',
625 => '1',
626 => '1',
627 => '0',
628 => '0',
629 => '0',
630 => '0',
631 => '0',
632 => '0',
633 => '0',
634 => '0',
635 => '0',
636 => '0',
637 => '0',
638 => '1',
639 => '1',
640 => '1',
641 => '1',
642 => '1',
643 => '0',
644 => '0',
645 => '0',
646 => '0',
647 => '0',
648 => '0',
649 => '0',
650 => '0',
651 => '0',
652 => '0',
653 => '0',
654 => '1',
655 => '1',
656 => '1',
657 => '1',
658 => '1',
659 => '0',
660 => '0',
661 => '0',
662 => '0',
663 => '0',
664 => '0',
665 => '0',
666 => '0',
667 => '0',
668 => '0',
669 => '0',
670 => '1',
671 => '1',
672 => '1',
673 => '1',
674 => '1',
675 => '0',
676 => '0',
677 => '0',
678 => '0',
679 => '0',
680 => '0',
681 => '0',
682 => '0',
683 => '0',
684 => '0',
685 => '0',
686 => '1',
687 => '1',
688 => '1',
689 => '1',
690 => '1',
691 => '0',
692 => '0',
693 => '0',
694 => '0',
695 => '0',
696 => '0',
697 => '0',
698 => '0',
699 => '0',
700 => '0',
701 => '0',
702 => '1',
703 => '1',
704 => '1',
705 => '1',
706 => '1',
707 => '0',
708 => '0',
709 => '0',
710 => '0',
711 => '0',
712 => '0',
713 => '0',
714 => '0',
715 => '0',
716 => '0',
717 => '0',
718 => '1',
719 => '1',
720 => '1',
721 => '1',
722 => '1',
723 => '0',
724 => '0',
725 => '0',
726 => '0',
727 => '0',
728 => '0',
729 => '0',
730 => '0',
731 => '0',
732 => '0',
733 => '0',
734 => '1',
735 => '1',
736 => '1',
737 => '1',
738 => '1',
739 => '0',
740 => '0',
741 => '0',
742 => '0',
743 => '0',
744 => '0',
745 => '0',
746 => '0',
747 => '0',
748 => '0',
749 => '0',
750 => '1',
751 => '1',
752 => '1',
753 => '1',
754 => '1',
755 => '0',
756 => '0',
757 => '0',
758 => '0',
759 => '0',
760 => '0',
761 => '0',
762 => '0',
763 => '0',
764 => '0',
765 => '0',
766 => '1',
767 => '1',
768 => '1',
769 => '1',
770 => '1',
771 => '0',
772 => '0',
773 => '0',
774 => '0',
775 => '0',
776 => '0',
777 => '0',
778 => '0',
779 => '0',
780 => '0',
781 => '0',
782 => '1',
783 => '1',
784 => '1',
785 => '1',
786 => '1',
787 => '0',
788 => '0',
789 => '0',
790 => '0',
791 => '0',
792 => '0',
793 => '0',
794 => '0',
795 => '0',
796 => '0',
797 => '0',
798 => '1',
799 => '1',
800 => '1',
801 => '1',
802 => '1',
803 => '0',
804 => '0',
805 => '0',
806 => '0',
807 => '0',
808 => '0',
809 => '0',
810 => '0',
811 => '0',
812 => '0',
813 => '0',
814 => '1',
815 => '1',
816 => '1',
817 => '1',
818 => '1',
819 => '0',
820 => '0',
821 => '0',
822 => '0',
823 => '0',
824 => '0',
825 => '0',
826 => '0',
827 => '0',
828 => '0',
829 => '0',
830 => '1',
831 => '1',
832 => '1',
833 => '1',
834 => '1',
835 => '0',
836 => '0',
837 => '0',
838 => '0',
839 => '0',
840 => '0',
841 => '0',
842 => '0',
843 => '0',
844 => '0',
845 => '0',
846 => '1',
847 => '1',
848 => '1',
849 => '1',
850 => '1',
851 => '0',
852 => '0',
853 => '0',
854 => '0',
855 => '0',
856 => '0',
857 => '0',
858 => '0',
859 => '0',
860 => '0',
861 => '0',
862 => '1',
863 => '1',
864 => '1',
865 => '1',
866 => '1',
867 => '0',
868 => '0',
869 => '0',
870 => '0',
871 => '0',
872 => '0',
873 => '0',
874 => '0',
875 => '0',
876 => '0',
877 => '0',
878 => '1',
879 => '1',
880 => '1',
881 => '1',
882 => '1',
883 => '0',
884 => '0',
885 => '0',
886 => '0',
887 => '0',
888 => '0',
889 => '0',
890 => '0',
891 => '0',
892 => '0',
893 => '0',
894 => '1',
895 => '1',
896 => '1',
897 => '1',
898 => '1',
899 => '0',
900 => '0',
901 => '0',
902 => '0',
903 => '0',
904 => '0',
905 => '0',
906 => '0',
907 => '0',
908 => '0',
909 => '0',
910 => '1',
911 => '1',
912 => '1',
913 => '1',
914 => '1',
915 => '0',
916 => '0',
917 => '0',
918 => '0',
919 => '0',
920 => '0',
921 => '0',
922 => '0',
923 => '0',
924 => '0',
925 => '0',
926 => '1',
927 => '1',
928 => '1',
929 => '1',
930 => '1',
931 => '0',
932 => '0',
933 => '0',
934 => '0',
935 => '0',
936 => '0',
937 => '0',
938 => '0',
939 => '0',
940 => '0',
941 => '0',
942 => '1',
943 => '1',
944 => '1',
945 => '1',
946 => '1',
947 => '0',
948 => '0',
949 => '0',
950 => '0',
951 => '0',
952 => '0',
953 => '0',
954 => '0',
955 => '0',
956 => '0',
957 => '0',
958 => '1',
959 => '1',
960 => '1',
961 => '1',
962 => '0',
963 => '0',
964 => '0',
965 => '0',
966 => '0',
967 => '0',
968 => '0',
969 => '0',
970 => '0',
971 => '0',
972 => '0',
973 => '1',
974 => '1',
975 => '1',
976 => '1',
977 => '1',
978 => '0',
979 => '0',
980 => '0',
981 => '0',
982 => '0',
983 => '0',
984 => '0',
985 => '0',
986 => '0',
987 => '0',
988 => '0',
989 => '1',
990 => '1',
991 => '1',
992 => '1',
993 => '1',
994 => '1',
995 => '1',
996 => '1',
997 => '0',
998 => '0',
999 => '0',
1000 => '0',
1001 => '0',
1002 => '0',
1003 => '0',
1004 => '1',
1005 => '1',
1006 => '1',
1007 => '1',
1008 => '1',
1009 => '1',
1010 => '1',
1011 => '1',
1012 => '1',
1013 => '1',
1014 => '0',
1015 => '0',
1016 => '0',
1017 => '0',
1018 => '0',
1019 => '1',
1020 => '1',
1021 => '1',
1022 => '1',
1023 => '1',
1024 => '1',
1025 => '1',
1026 => '1',
1027 => '1',
1028 => '1',
1029 => '1',
1030 => '1',
1031 => '1',
1032 => '1',
1033 => '1',
1034 => '1',
1035 => '1',
1036 => '1',
1037 => '1',
1038 => '1',
1039 => '1',
1040 => '1',
1041 => '1',
1042 => '1',
1043 => '0',
1044 => '0',
1045 => '0',
1046 => '1',
1047 => '1',
1048 => '1',
1049 => '1',
1050 => '1',
1051 => '1',
1052 => '1',
1053 => '1',
1054 => '1',
1055 => '1',
1056 => '1',
1057 => '1',
1058 => '0',
1059 => '0',
1060 => '0',
1061 => '0',
1062 => '0',
1063 => '1',
1064 => '1',
1065 => '1',
1066 => '1',
1067 => '1',
1068 => '1',
1069 => '1',
1070 => '1',
1071 => '1',
1072 => '1',
1073 => '0',
1074 => '0',
1075 => '0',
1076 => '0',
1077 => '0',
1078 => '0',
1079 => '0',
1080 => '0',
1081 => '1',
1082 => '1',
1083 => '1',
1084 => '1',
1085 => '1',
1086 => '1',
1087 => '1',
1088 => '0',
1089 => '0',
1090 => '0',
1091 => '0',
1092 => '0',
1093 => '0',
1094 => '0',
1095 => '0',
1096 => '0',
1097 => '0',
1098 => '1',
1099 => '1',
1100 => '1',
1101 => '1',
1102 => '1',
1103 => '1',
1104 => '0',
1105 => '0',
1106 => '0',
1107 => '0',
1108 => '0',
1109 => '0',
1110 => '0',
1111 => '0',
1112 => '0',
1113 => '0',
1114 => '0',
1115 => '0',
1116 => '1',
1117 => '1',
1118 => '1',
1119 => '1',
1120 => '0',
1121 => '0',
1122 => '0',
1123 => '0',
1124 => '0',
1125 => '0',
1126 => '0',
1127 => '0',
1128 => '0',
1129 => '0',
1130 => '0',
1131 => '0',
1132 => '0',
1133 => '1',
1134 => '1',
1135 => '1',
1136 => '1',
1137 => '0',
1138 => '0',
1139 => '0',
1140 => '0',
1141 => '0',
1142 => '0',
1143 => '0',
1144 => '0',
1145 => '0',
1146 => '0',
1147 => '0',
1148 => '0',
1149 => '0',
1150 => '1',
1151 => '1',
1152 => '1',
1153 => '1',
1154 => '0',
1155 => '0',
1156 => '0',
1157 => '0',
1158 => '0',
1159 => '0',
1160 => '0',
1161 => '0',
1162 => '0',
1163 => '0',
1164 => '0',
1165 => '0',
1166 => '0',
1167 => '1',
1168 => '1',
1169 => '1',
1170 => '1',
1171 => '0',
1172 => '0',
1173 => '0',
1174 => '0',
1175 => '0',
1176 => '0',
1177 => '0',
1178 => '0',
1179 => '0',
1180 => '0',
1181 => '0',
1182 => '0',
1183 => '0',
1184 => '1',
1185 => '1',
1186 => '1',
1187 => '1',
1188 => '0',
1189 => '0',
1190 => '0',
1191 => '0',
1192 => '0',
1193 => '0',
1194 => '0',
1195 => '0',
1196 => '0',
1197 => '0',
1198 => '0',
1199 => '0',
1200 => '1',
1201 => '1',
1202 => '1',
1203 => '1',
1204 => '1',
1205 => '0',
1206 => '0',
1207 => '0',
1208 => '0',
1209 => '0',
1210 => '0',
1211 => '0',
1212 => '0',
1213 => '0',
1214 => '0',
1215 => '0',
1216 => '1',
1217 => '1',
1218 => '1',
1219 => '1',
1220 => '1',
1221 => '1',
1222 => '0',
1223 => '0',
1224 => '0',
1225 => '0',
1226 => '0',
1227 => '0',
1228 => '0',
1229 => '0',
1230 => '0',
1231 => '1',
1232 => '1',
1233 => '1',
1234 => '1',
1235 => '1',
1236 => '1',
1237 => '1',
1238 => '1',
1239 => '0',
1240 => '0',
1241 => '0',
1242 => '0',
1243 => '0',
1244 => '0',
1245 => '0',
1246 => '0',
1247 => '1',
1248 => '1',
1249 => '1',
1250 => '1',
1251 => '1',
1252 => '1',
1253 => '1',
1254 => '1',
1255 => '1',
1256 => '1',
1257 => '0',
1258 => '0',
1259 => '0',
1260 => '0',
1261 => '0',
1262 => '1',
1263 => '1',
1264 => '1',
1265 => '1',
1266 => '1',
1267 => '1',
1268 => '1',
1269 => '1',
1270 => '1',
1271 => '1',
1272 => '1',
1273 => '1',
1274 => '1',
1275 => '0',
1276 => '0',
1277 => '1',
1278 => '1',
1279 => '1',
1280 => '1',
1281 => '1',
1282 => '1',
1283 => '1',
1284 => '1',
1285 => '1',
1286 => '1',
1287 => '1',
1288 => '1',
1289 => '1',
1290 => '1',
1291 => '1',
1292 => '1',
1293 => '1',
1294 => '1',
1295 => '1',
1296 => '1',
1297 => '1',
1298 => '1',
1299 => '1',
1300 => '1',
1301 => '0',
1302 => '0',
1303 => '0',
1304 => '0',
1305 => '0',
1306 => '0',
1307 => '1',
1308 => '1',
1309 => '1',
1310 => '1',
1311 => '1',
1312 => '1',
1313 => '1',
1314 => '1',
1315 => '1',
1316 => '0',
1317 => '0',
1318 => '0',
1319 => '0',
1320 => '0',
1321 => '0',
1322 => '0',
1323 => '0',
1324 => '1',
1325 => '1',
1326 => '1',
1327 => '1',
1328 => '1',
1329 => '1',
1330 => '1',
1331 => '0',
1332 => '0',
1333 => '0',
1334 => '0',
1335 => '0',
1336 => '0',
1337 => '0',
1338 => '0',
1339 => '0',
1340 => '0',
1341 => '1',
1342 => '1',
1343 => '1',
1344 => '1',
1345 => '1',
1346 => '1',
1347 => '0',
1348 => '0',
1349 => '0',
1350 => '0',
1351 => '0',
1352 => '0',
1353 => '0',
1354 => '0',
1355 => '0',
1356 => '0',
1357 => '1',
1358 => '1',
1359 => '1',
1360 => '1',
1361 => '1',
1362 => '1',
1363 => '0',
1364 => '0',
1365 => '0',
1366 => '0',
1367 => '0',
1368 => '0',
1369 => '0',
1370 => '0',
1371 => '0',
1372 => '0',
1373 => '1',
1374 => '1',
1375 => '1',
1376 => '1',
1377 => '1',
1378 => '1',
1379 => '0',
1380 => '0',
1381 => '0',
1382 => '0',
1383 => '0',
1384 => '0',
1385 => '0',
1386 => '0',
1387 => '0',
1388 => '0',
1389 => '1',
1390 => '1',
1391 => '1',
1392 => '1',
1393 => '1',
1394 => '1',
1395 => '0',
1396 => '0',
1397 => '0',
1398 => '0',
1399 => '0',
1400 => '0',
1401 => '0',
1402 => '0',
1403 => '0',
1404 => '0',
1405 => '1',
1406 => '1',
1407 => '1',
1408 => '1',
1409 => '1',
1410 => '1',
1411 => '0',
1412 => '0',
1413 => '0',
1414 => '0',
1415 => '0',
1416 => '0',
1417 => '0',
1418 => '0',
1419 => '0',
1420 => '0',
1421 => '1',
1422 => '1',
1423 => '1',
1424 => '1',
1425 => '1',
1426 => '1',
1427 => '0',
1428 => '0',
1429 => '0',
1430 => '0',
1431 => '0',
1432 => '0',
1433 => '0',
1434 => '0',
1435 => '0',
1436 => '0',
1437 => '1',
1438 => '1',
1439 => '1',
1440 => '1',
1441 => '1',
1442 => '1',
1443 => '0',
1444 => '0',
1445 => '0',
1446 => '0',
1447 => '0',
1448 => '0',
1449 => '0',
1450 => '0',
1451 => '0',
1452 => '0',
1453 => '1',
1454 => '1',
1455 => '1',
1456 => '1',
1457 => '1',
1458 => '1',
1459 => '0',
1460 => '0',
1461 => '0',
1462 => '0',
1463 => '0',
1464 => '0',
1465 => '0',
1466 => '0',
1467 => '0',
1468 => '0',
1469 => '1',
1470 => '1',
1471 => '1',
1472 => '1',
1473 => '1',
1474 => '1',
1475 => '0',
1476 => '0',
1477 => '0',
1478 => '0',
1479 => '0',
1480 => '0',
1481 => '0',
1482 => '0',
1483 => '0',
1484 => '0',
1485 => '1',
1486 => '1',
1487 => '1',
1488 => '1',
1489 => '1',
1490 => '1',
1491 => '1',
1492 => '0',
1493 => '0',
1494 => '0',
1495 => '0',
1496 => '0',
1497 => '0',
1498 => '0',
1499 => '0',
1500 => '1',
1501 => '1',
1502 => '1',
1503 => '1',
1504 => '1',
1505 => '1',
1506 => '1',
1507 => '1',
1508 => '1',
1509 => '0',
1510 => '0',
1511 => '0',
1512 => '0',
1513 => '0',
1514 => '0',
1515 => '1',
1516 => '1',
1517 => '1',
1518 => '1',
1519 => '1',
1520 => '1',
1521 => '1',
1522 => '1',
1523 => '1',
1524 => '1',
1525 => '1',
1526 => '1',
1527 => '1',
1528 => '1',
1529 => '1',
1530 => '1',
1531 => '1',
1532 => '1',
1533 => '1',
1534 => '1',
1535 => '1',
1536 => '1',
1537 => '1',
1538 => '1',
1539 => '1',
1540 => '1',
1541 => '1',
1542 => '1',
1543 => '1',
1544 => '1',
1545 => '1',
1546 => '1',
1547 => '1',
1548 => '1',
1549 => '1',
1550 => '1',
1551 => '1',
1552 => '1',
1553 => '1',
1554 => '1',
1555 => '1',
1556 => '1',
1557 => '1',
1558 => '1',
1559 => '1',
1560 => '1',
1561 => '1',
1562 => '1',
1563 => '0',
1564 => '0',
1565 => '1',
1566 => '1',
1567 => '1',
1568 => '1',
1569 => '1',
1570 => '1',
1571 => '1',
1572 => '1',
1573 => '1',
1574 => '1',
1575 => '1',
1576 => '1',
1577 => '1',
1578 => '0',
1579 => '0',
1580 => '0',
1581 => '0',
1582 => '1',
1583 => '1',
1584 => '1',
1585 => '1',
1586 => '1',
1587 => '1',
1588 => '1',
1589 => '1',
1590 => '1',
1591 => '1',
1592 => '0',
1593 => '0',
1594 => '0',
1595 => '0',
1596 => '0',
1597 => '0',
1598 => '0',
1599 => '1',
1600 => '1',
1601 => '1',
1602 => '1',
1603 => '1',
1604 => '1',
1605 => '1',
1606 => '0',
1607 => '0',
1608 => '0',
1609 => '0',
1610 => '0',
1611 => '0',
1612 => '0',
1613 => '0',
1614 => '0',
1615 => '0',
1616 => '1',
1617 => '1',
1618 => '1',
1619 => '1',
1620 => '1',
1621 => '0',
1622 => '0',
1623 => '0',
1624 => '0',
1625 => '0',
1626 => '0',
1627 => '0',
1628 => '0',
1629 => '0',
1630 => '0',
1631 => '0',
1632 => '1',
1633 => '1',
1634 => '1',
1635 => '0',
1636 => '0',
1637 => '0',
1638 => '0',
1639 => '0',
1640 => '0',
1641 => '0',
1642 => '0',
1643 => '0',
1644 => '0',
1645 => '0',
1646 => '0',
1647 => '0',
1648 => '1',
1649 => '1',
1650 => '0',
1651 => '0',
1652 => '0',
1653 => '0',
1654 => '0',
1655 => '0',
1656 => '0',
1657 => '0',
1658 => '0',
1659 => '0',
1660 => '0',
1661 => '0',
1662 => '0',
1663 => '0',
1664 => '1',
1665 => '0',
1666 => '0',
1667 => '0',
1668 => '0',
1669 => '0',
1670 => '0',
1671 => '0',
1672 => '0',
1673 => '0',
1674 => '0',
1675 => '0',
1676 => '0',
1677 => '0',
1678 => '0',
1679 => '1',
1680 => '0',
1681 => '0',
1682 => '0',
1683 => '0',
1684 => '0',
1685 => '0',
1686 => '0',
1687 => '0',
1688 => '0',
1689 => '0',
1690 => '0',
1691 => '0',
1692 => '0',
1693 => '0',
1694 => '1',
1695 => '1',
1696 => '0',
1697 => '0',
1698 => '0',
1699 => '0',
1700 => '0',
1701 => '0',
1702 => '0',
1703 => '0',
1704 => '0',
1705 => '0',
1706 => '0',
1707 => '0',
1708 => '0',
1709 => '1',
1710 => '1',
1711 => '1',
1712 => '0',
1713 => '0',
1714 => '0',
1715 => '0',
1716 => '0',
1717 => '0',
1718 => '0',
1719 => '0',
1720 => '0',
1721 => '0',
1722 => '0',
1723 => '0',
1724 => '1',
1725 => '1',
1726 => '1',
1727 => '1',
1728 => '1',
1729 => '0',
1730 => '0',
1731 => '0',
1732 => '0',
1733 => '0',
1734 => '0',
1735 => '0',
1736 => '0',
1737 => '0',
1738 => '1',
1739 => '1',
1740 => '1',
1741 => '1',
1742 => '1',
1743 => '1',
1744 => '1',
1745 => '1',
1746 => '0',
1747 => '0',
1748 => '0',
1749 => '0',
1750 => '0',
1751 => '0',
1752 => '0',
1753 => '1',
1754 => '1',
1755 => '1',
1756 => '1',
1757 => '1',
1758 => '1',
1759 => '1',
1760 => '1',
1761 => '1',
1762 => '1',
1763 => '0',
1764 => '0',
1765 => '0',
1766 => '0',
1767 => '0',
1768 => '1',
1769 => '1',
1770 => '1',
1771 => '1',
1772 => '1',
1773 => '1',
1774 => '1',
1775 => '1',
1776 => '1',
1777 => '1',
1778 => '1',
1779 => '1',
1780 => '0',
1781 => '0',
1782 => '1',
1783 => '1',
1784 => '1',
1785 => '1',
1786 => '1',
1787 => '1',
1788 => '1',
1789 => '1',
1790 => '1',
1791 => '1',
1792 => '1',
1793 => '1',
1794 => '1',
1795 => '1',
1796 => '1',
1797 => '1',
1798 => '1',
1799 => '1',
1800 => '1',
1801 => '1',
1802 => '1',
1803 => '1',
1804 => '1',
1805 => '1',
1806 => '1',
1807 => '1',
1808 => '1',
1809 => '1',
1810 => '1',
1811 => '1',
1812 => '1',
1813 => '1',
1814 => '1',
1815 => '1',
1816 => '1',
1817 => '1',
1818 => '1',
1819 => '1',
1820 => '1',
1821 => '1',
1822 => '1',
1823 => '1',
1824 => '1',
1825 => '1',
1826 => '1',
1827 => '1',
1828 => '1',
1829 => '1',
1830 => '1',
1831 => '1',
1832 => '1',
1833 => '1',
1834 => '1',
1835 => '1',
1836 => '1',
1837 => '1',
1838 => '1',
1839 => '1',
1840 => '1',
1841 => '1',
1842 => '0',
1843 => '0',
1844 => '0',
1845 => '0',
1846 => '0',
1847 => '0',
1848 => '0',
1849 => '0',
1850 => '0',
1851 => '0',
1852 => '0',
1853 => '0',
1854 => '1',
1855 => '1',
1856 => '1',
1857 => '0',
1858 => '0',
1859 => '0',
1860 => '0',
1861 => '0',
1862 => '0',
1863 => '0',
1864 => '0',
1865 => '0',
1866 => '0',
1867 => '0',
1868 => '0',
1869 => '0',
1870 => '0',
1871 => '1',
1872 => '0',
1873 => '0',
1874 => '0',
1875 => '0',
1876 => '0',
1877 => '0',
1878 => '0',
1879 => '0',
1880 => '0',
1881 => '0',
1882 => '0',
1883 => '0',
1884 => '0',
1885 => '0',
1886 => '0',
1887 => '0',
1888 => '0',
1889 => '0',
1890 => '0',
1891 => '0',
1892 => '0',
1893 => '0',
1894 => '0',
1895 => '0',
1896 => '0',
1897 => '0',
1898 => '0',
1899 => '0',
1900 => '0',
1901 => '0',
1902 => '0',
1903 => '0',
1904 => '0',
1905 => '0',
1906 => '0',
1907 => '0',
1908 => '0',
1909 => '0',
1910 => '0',
1911 => '0',
1912 => '0',
1913 => '0',
1914 => '0',
1915 => '0',
1916 => '0',
1917 => '0',
1918 => '0',
1919 => '0',
1920 => '0',
1921 => '0',
1922 => '0',
1923 => '0',
1924 => '0',
1925 => '0',
1926 => '0',
1927 => '0',
1928 => '0',
1929 => '0',
1930 => '0',
1931 => '0',
1932 => '0',
1933 => '0',
1934 => '0',
1935 => '0',
1936 => '0',
1937 => '0',
1938 => '0',
1939 => '0',
1940 => '0',
1941 => '0',
1942 => '0',
1943 => '0',
1944 => '0',
1945 => '0',
1946 => '0',
1947 => '0',
1948 => '0',
1949 => '0',
1950 => '0',
1951 => '0',
1952 => '0',
1953 => '0',
1954 => '0',
1955 => '0',
1956 => '0',
1957 => '0',
1958 => '0',
1959 => '0',
1960 => '0',
1961 => '0',
1962 => '0',
1963 => '0',
1964 => '0',
1965 => '0',
1966 => '0',
1967 => '0',
1968 => '1',
1969 => '0',
1970 => '0',
1971 => '0',
1972 => '0',
1973 => '0',
1974 => '0',
1975 => '0',
1976 => '0',
1977 => '0',
1978 => '0',
1979 => '0',
1980 => '0',
1981 => '0',
1982 => '0',
1983 => '1',
1984 => '1',
1985 => '1',
1986 => '0',
1987 => '0',
1988 => '0',
1989 => '0',
1990 => '0',
1991 => '0',
1992 => '0',
1993 => '0',
1994 => '0',
1995 => '0',
1996 => '0',
1997 => '0',
1998 => '1',
1999 => '1',
2000 => '1',
2001 => '1',
2002 => '1',
2003 => '1',
2004 => '1',
2005 => '1',
2006 => '1',
2007 => '1',
2008 => '1',
2009 => '1',
2010 => '1',
2011 => '1',
2012 => '1',
2013 => '1',
2014 => '1',
2015 => '1',
2016 => '1',
2017 => '1',
2018 => '1',
2019 => '1',
2020 => '1',
2021 => '1',
2022 => '1',
2023 => '1',
2024 => '1',
2025 => '1',
2026 => '1',
2027 => '1',
2028 => '1',
2029 => '1',
2030 => '1',
2031 => '1',
2032 => '1',
2033 => '1',
2034 => '1',
2035 => '1',
2036 => '1',
2037 => '1',
2038 => '1',
2039 => '1',
2040 => '1',
2041 => '1',
2042 => '1',
2043 => '1',
2044 => '1',
2045 => '1',
2046 => '1',
2047 => '1',
        others => '1'
    );
begin
 
    -- G?n?ration: d?tection de collision pixel / acteur
    gen_actor_check: for i in 0 to 7 generate
    begin
        s_actor_hit(i) <= '1' when (
            to_integer(unsigned(i_view_x)) >= to_integer(unsigned(actor_pos_x(i))) and
            to_integer(unsigned(i_view_x)) <  to_integer(unsigned(actor_pos_x(i))) + 16 and
            to_integer(unsigned(i_view_y)) >= to_integer(unsigned(actor_pos_y(i))) and
            to_integer(unsigned(i_view_y)) <  to_integer(unsigned(actor_pos_y(i))) + 16
        ) else '0';
    end generate;
    
    process(i_clk)
      variable writeIndex : std_logic_vector (11 downto 0);
      variable writeIndex_int : integer;
      variable writeData : std_logic;
      begin
        if rising_edge(i_clk) then
            if i_ch_we = '1' then
                writeIndex := i_tile_id_write & i_ch_y & i_ch_x;
                writeIndex_int := to_integer(unsigned(writeIndex));
                writeData := '0';
                if i_ch_cc = "1111" then
                    writeData := '1';
                end if;
                tile_data_map_a(writeIndex_int) <= writeData;
            end if;
        end if;
      end process;
 
    -- R�solution: acteur de plus haute priorit� (ID plus bas)
    process(i_clk)
        variable rel_x, rel_y : integer range 0 to 15;
        variable pix_x_flipped : std_logic_vector (3 downto 0);
        variable pix_y_flipped : std_logic_vector (3 downto 0);
        variable index : std_logic_vector (11 downto 0);
        variable index_int : integer;
        variable pix_x : std_logic_vector (3 downto 0);
        variable pix_y : std_logic_vector (3 downto 0);
        variable pix_x_int : integer;
        variable pix_y_int : integer;
        variable flip_x : std_logic;
        variable flip_y : std_logic;
        variable tileId : std_logic_vector (3 downto 0);
    begin
    if rising_edge(i_clk) then
        -- Default values
        o_tile_id <= (others => '0');
        o_flip_x <= '0';
        o_flip_y <= '0';
        o_pix_x <= (others => '0');
        o_pix_y <= (others => '0');
        o_is_actor_present <= '0';
        -- Priority loop: lowest i with hit gets selected and non transparent
        for i in 0 to 7 loop
            if s_actor_hit(i) = '1' then
                rel_x := to_integer(unsigned(i_view_x)) - to_integer(unsigned(actor_pos_x(i)));
                rel_y := to_integer(unsigned(i_view_y)) - to_integer(unsigned(actor_pos_y(i)));
                pix_x := std_logic_vector(to_unsigned(rel_x, 4));
                pix_y := std_logic_vector(to_unsigned(rel_y, 4));
                flip_x := actor_flip_x(i);
                flip_y := actor_flip_y(i);
                tileId := actor_tile_id(i);
                pix_x_int := to_integer(unsigned(pix_x));
                pix_y_int := to_integer(unsigned(pix_y));
                if flip_x = '1' then
                    pix_x_flipped := std_logic_vector(to_unsigned(15 - pix_x_int, 4));
                else
                    pix_x_flipped := pix_x;
                end if;
                if flip_y = '1' then
                    pix_y_flipped := std_logic_vector(to_unsigned(15 - pix_y_int, 4));
                else
                    pix_y_flipped := pix_y;
                end if;
                index := tileId & pix_y_flipped & pix_x_flipped;
                index_int := to_integer(unsigned(index));
            
                if tile_data_map_a(index_int) = '0' then
                    o_tile_id <= tileId;
                    o_flip_x <= flip_x;
                    o_flip_y <= flip_y;
                    o_pix_x <= pix_x;
                    o_pix_y <= pix_y;
                    o_is_actor_present <= '1';
                end if;
            end if;
        end loop;
        end if;
    end process;
    -- ?criture des donn?es d'acteurs
    process(i_clk)
        variable id : integer;
    begin
        if rising_edge(i_clk) then
            id := to_integer(unsigned(i_act_id));
 
            if i_ch_setpos = '1' then
                actor_pos_x(id) <= i_newpos_x;
                actor_pos_y(id) <= i_newpos_y;
            end if;
 
            if i_ch_tile_id = '1' then
                actor_tile_id(id) <= i_tile_id;
            end if;
 
            if i_ch_flipX = '1' then
                actor_flip_x(id) <= i_flip_x;
            end if;
 
            if i_ch_flipY = '1' then
                actor_flip_y(id) <= i_flip_y;
            end if;
        end if;
    end process;
 
end Behavioral;
