library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity TuileBackBuff2 is
    Port(
    i_x : in STD_LOGIC_VECTOR (2 downto 0);
    i_y : in STD_LOGIC_VECTOR (2 downto 0);
    i_tile_id : in STD_LOGIC_VECTOR (4 downto 0);
    i_ch_x : in STD_LOGIC_VECTOR (2 downto 0);
    i_ch_y : in STD_LOGIC_VECTOR (2 downto 0);
    i_ch_cc : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_we : in std_logic;
    i_clk : in STD_LOGIC;
    i_flip_y : in STD_LOGIC;
    i_tile_id_write : in STD_LOGIC_VECTOR (4 downto 0);
    o_colorCode : out STD_LOGIC_VECTOR (3 downto 0));
end TuileBackBuff2;

architecture Behavioral of TuileBackBuff2 is
constant wh : std_logic_vector (3 downto 0) := "0000"; -- White
constant bl : std_logic_vector (3 downto 0) := "0001"; -- Black
constant ye : std_logic_vector (3 downto 0) := "0010"; -- Yellow
constant dg : std_logic_vector (3 downto 0) := "0011"; -- Dark Green
constant oa : std_logic_vector (3 downto 0) := "0100"; -- Orange
constant bu : std_logic_vector (3 downto 0) := "0101"; -- Blue
constant ge : std_logic_vector (3 downto 0) := "0110"; -- Green
constant lo : std_logic_vector (3 downto 0) := "0111"; -- Light Brown
constant br : std_logic_vector (3 downto 0) := "1000"; -- Brown
constant lg : std_logic_vector (3 downto 0) := "1001"; -- Light Gray
constant gr : std_logic_vector (3 downto 0) := "1010"; -- Gray
constant lb : std_logic_vector (3 downto 0) := "1011"; -- Light Blue
constant sb : std_logic_vector (3 downto 0) := "1100"; -- Sky Blue
constant sa : std_logic_vector (3 downto 0) := "1101"; -- Salmon
constant pi : std_logic_vector (3 downto 0) := "1110"; -- Pink
constant pu : std_logic_vector (3 downto 0) := "1111"; -- Purple
    
    type tile_d_array_t is array (0 to 2047) of std_logic_vector(3 downto 0);
    signal tile_data_map_d : tile_d_array_t :=
    (
        0 => wh,
1 => wh,
2 => wh,
3 => wh,
4 => wh,
5 => wh,
6 => wh,
7 => wh,
8 => wh,
9 => wh,
10 => wh,
11 => wh,
12 => wh,
13 => wh,
14 => wh,
15 => wh,
16 => wh,
17 => wh,
18 => wh,
19 => wh,
20 => wh,
21 => wh,
22 => wh,
23 => wh,
24 => wh,
25 => wh,
26 => wh,
27 => wh,
28 => wh,
29 => wh,
30 => wh,
31 => wh,
32 => wh,
33 => wh,
34 => wh,
35 => wh,
36 => wh,
37 => wh,
38 => wh,
39 => wh,
40 => wh,
41 => wh,
42 => wh,
43 => wh,
44 => wh,
45 => wh,
46 => wh,
47 => wh,
48 => wh,
49 => wh,
50 => wh,
51 => wh,
52 => wh,
53 => wh,
54 => wh,
55 => wh,
56 => wh,
57 => wh,
58 => wh,
59 => wh,
60 => wh,
61 => wh,
62 => wh,
63 => wh,
64 => wh,
65 => wh,
66 => sb,
67 => lb,
68 => lb,
69 => sb,
70 => wh,
71 => wh,
72 => wh,
73 => wh,
74 => sb,
75 => lb,
76 => lb,
77 => sb,
78 => sb,
79 => wh,
80 => wh,
81 => wh,
82 => sb,
83 => lb,
84 => lb,
85 => sb,
86 => wh,
87 => wh,
88 => wh,
89 => sb,
90 => lb,
91 => lb,
92 => lb,
93 => sb,
94 => wh,
95 => wh,
96 => wh,
97 => wh,
98 => sb,
99 => lb,
100 => lb,
101 => sb,
102 => wh,
103 => wh,
104 => wh,
105 => wh,
106 => sb,
107 => lb,
108 => lb,
109 => sb,
110 => sb,
111 => wh,
112 => wh,
113 => sb,
114 => sb,
115 => lb,
116 => lb,
117 => sb,
118 => wh,
119 => wh,
120 => wh,
121 => wh,
122 => sb,
123 => lb,
124 => lb,
125 => sb,
126 => wh,
127 => wh,
128 => wh,
129 => wh,
130 => pi,
131 => sa,
132 => sa,
133 => pi,
134 => wh,
135 => wh,
136 => wh,
137 => wh,
138 => pi,
139 => sa,
140 => sa,
141 => pi,
142 => wh,
143 => wh,
144 => wh,
145 => pi,
146 => pi,
147 => sa,
148 => sa,
149 => pi,
150 => wh,
151 => wh,
152 => wh,
153 => wh,
154 => pi,
155 => sa,
156 => sa,
157 => pi,
158 => wh,
159 => wh,
160 => wh,
161 => wh,
162 => pi,
163 => sa,
164 => sa,
165 => sa,
166 => pi,
167 => wh,
168 => wh,
169 => wh,
170 => pi,
171 => sa,
172 => sa,
173 => pi,
174 => wh,
175 => wh,
176 => wh,
177 => pi,
178 => pi,
179 => sa,
180 => sa,
181 => pi,
182 => wh,
183 => wh,
184 => wh,
185 => wh,
186 => pi,
187 => sa,
188 => sa,
189 => pi,
190 => wh,
191 => wh,
192 => wh,
193 => wh,
194 => wh,
195 => wh,
196 => wh,
197 => wh,
198 => wh,
199 => wh,
200 => wh,
201 => wh,
202 => wh,
203 => wh,
204 => wh,
205 => lg,
206 => lg,
207 => pi,
208 => wh,
209 => wh,
210 => wh,
211 => lg,
212 => lg,
213 => lg,
214 => lg,
215 => wh,
216 => wh,
217 => wh,
218 => lg,
219 => lg,
220 => lg,
221 => wh,
222 => gr,
223 => lg,
224 => wh,
225 => wh,
226 => lg,
227 => lg,
228 => gr,
229 => lg,
230 => lg,
231 => lg,
232 => wh,
233 => lg,
234 => wh,
235 => gr,
236 => wh,
237 => gr,
238 => lg,
239 => lg,
240 => wh,
241 => wh,
242 => wh,
243 => wh,
244 => lg,
245 => gr,
246 => lg,
247 => wh,
248 => wh,
249 => wh,
250 => wh,
251 => wh,
252 => wh,
253 => wh,
254 => wh,
255 => lg,
256 => lg,
257 => lg,
258 => wh,
259 => lg,
260 => lg,
261 => lg,
262 => lg,
263 => wh,
264 => wh,
265 => wh,
266 => wh,
267 => pi,
268 => wh,
269 => pi,
270 => wh,
271 => lg,
272 => wh,
273 => pi,
274 => wh,
275 => pi,
276 => pi,
277 => wh,
278 => pi,
279 => pi,
280 => lg,
281 => wh,
282 => lg,
283 => pi,
284 => gr,
285 => pi,
286 => lg,
287 => gr,
288 => pi,
289 => lg,
290 => lg,
291 => gr,
292 => gr,
293 => gr,
294 => gr,
295 => lg,
296 => gr,
297 => gr,
298 => gr,
299 => lg,
300 => gr,
301 => gr,
302 => lg,
303 => gr,
304 => wh,
305 => gr,
306 => gr,
307 => gr,
308 => pi,
309 => gr,
310 => gr,
311 => gr,
312 => wh,
313 => wh,
314 => wh,
315 => wh,
316 => gr,
317 => wh,
318 => gr,
319 => pi,
320 => wh,
321 => wh,
322 => wh,
323 => wh,
324 => wh,
325 => wh,
326 => wh,
327 => wh,
328 => lg,
329 => lg,
330 => wh,
331 => wh,
332 => wh,
333 => wh,
334 => wh,
335 => wh,
336 => gr,
337 => gr,
338 => gr,
339 => gr,
340 => wh,
341 => wh,
342 => wh,
343 => wh,
344 => pi,
345 => pi,
346 => lg,
347 => gr,
348 => gr,
349 => wh,
350 => wh,
351 => wh,
352 => pi,
353 => gr,
354 => gr,
355 => lg,
356 => lg,
357 => wh,
358 => wh,
359 => wh,
360 => gr,
361 => lg,
362 => gr,
363 => gr,
364 => lg,
365 => gr,
366 => wh,
367 => wh,
368 => gr,
369 => gr,
370 => pi,
371 => lg,
372 => pi,
373 => gr,
374 => wh,
375 => wh,
376 => gr,
377 => pi,
378 => pi,
379 => wh,
380 => wh,
381 => pi,
382 => wh,
383 => wh,
384 => wh,
385 => wh,
386 => wh,
387 => wh,
388 => wh,
389 => wh,
390 => wh,
391 => wh,
392 => wh,
393 => wh,
394 => wh,
395 => pi,
396 => lg,
397 => pi,
398 => lg,
399 => wh,
400 => wh,
401 => wh,
402 => pi,
403 => wh,
404 => lg,
405 => pi,
406 => wh,
407 => pi,
408 => wh,
409 => pi,
410 => lg,
411 => pi,
412 => lg,
413 => lg,
414 => lg,
415 => wh,
416 => wh,
417 => lg,
418 => wh,
419 => lg,
420 => lg,
421 => lg,
422 => lg,
423 => lg,
424 => lg,
425 => lg,
426 => lg,
427 => pi,
428 => lg,
429 => lg,
430 => wh,
431 => lg,
432 => wh,
433 => lg,
434 => pi,
435 => lg,
436 => gr,
437 => pi,
438 => lg,
439 => gr,
440 => lg,
441 => lg,
442 => lg,
443 => lg,
444 => lg,
445 => lg,
446 => gr,
447 => gr,
448 => lg,
449 => wh,
450 => lg,
451 => lg,
452 => pi,
453 => gr,
454 => gr,
455 => gr,
456 => wh,
457 => pi,
458 => gr,
459 => lg,
460 => gr,
461 => lg,
462 => gr,
463 => gr,
464 => lg,
465 => lg,
466 => lg,
467 => gr,
468 => gr,
469 => gr,
470 => lg,
471 => pi,
472 => lg,
473 => gr,
474 => gr,
475 => gr,
476 => gr,
477 => lg,
478 => gr,
479 => lg,
480 => lg,
481 => pi,
482 => gr,
483 => gr,
484 => gr,
485 => gr,
486 => lg,
487 => gr,
488 => lg,
489 => pi,
490 => gr,
491 => gr,
492 => lg,
493 => lg,
494 => gr,
495 => lg,
496 => wh,
497 => gr,
498 => wh,
499 => lg,
500 => gr,
501 => pi,
502 => gr,
503 => pi,
504 => wh,
505 => wh,
506 => gr,
507 => wh,
508 => wh,
509 => gr,
510 => wh,
511 => wh,
512 => pi,
513 => wh,
514 => pi,
515 => pi,
516 => pi,
517 => gr,
518 => wh,
519 => wh,
520 => lg,
521 => gr,
522 => pi,
523 => lg,
524 => gr,
525 => gr,
526 => gr,
527 => wh,
528 => gr,
529 => gr,
530 => gr,
531 => gr,
532 => gr,
533 => gr,
534 => gr,
535 => gr,
536 => lg,
537 => gr,
538 => lg,
539 => gr,
540 => gr,
541 => gr,
542 => gr,
543 => wh,
544 => lg,
545 => gr,
546 => gr,
547 => gr,
548 => lg,
549 => gr,
550 => wh,
551 => gr,
552 => gr,
553 => gr,
554 => gr,
555 => gr,
556 => gr,
557 => gr,
558 => gr,
559 => wh,
560 => wh,
561 => gr,
562 => lg,
563 => gr,
564 => pi,
565 => pi,
566 => pi,
567 => gr,
568 => wh,
569 => pi,
570 => wh,
571 => pi,
572 => pi,
573 => wh,
574 => wh,
575 => pi,
576 => wh,
577 => wh,
578 => sb,
579 => lb,
580 => lb,
581 => sb,
582 => wh,
583 => wh,
584 => wh,
585 => wh,
586 => sb,
587 => sb,
588 => lb,
589 => sb,
590 => wh,
591 => wh,
592 => wh,
593 => wh,
594 => wh,
595 => lb,
596 => lb,
597 => wh,
598 => wh,
599 => wh,
600 => wh,
601 => wh,
602 => wh,
603 => sb,
604 => lb,
605 => wh,
606 => wh,
607 => wh,
608 => wh,
609 => wh,
610 => sb,
611 => wh,
612 => sb,
613 => wh,
614 => wh,
615 => wh,
616 => wh,
617 => wh,
618 => wh,
619 => lb,
620 => sb,
621 => wh,
622 => wh,
623 => wh,
624 => wh,
625 => wh,
626 => wh,
627 => sb,
628 => wh,
629 => wh,
630 => wh,
631 => wh,
632 => wh,
633 => wh,
634 => wh,
635 => wh,
636 => wh,
637 => wh,
638 => wh,
639 => wh,
640 => wh,
641 => wh,
642 => pi,
643 => sa,
644 => pi,
645 => pi,
646 => wh,
647 => wh,
648 => wh,
649 => wh,
650 => pi,
651 => sa,
652 => sa,
653 => pi,
654 => wh,
655 => wh,
656 => wh,
657 => wh,
658 => pi,
659 => pi,
660 => sa,
661 => pi,
662 => wh,
663 => wh,
664 => wh,
665 => wh,
666 => wh,
667 => sa,
668 => pi,
669 => wh,
670 => wh,
671 => wh,
672 => wh,
673 => wh,
674 => wh,
675 => pi,
676 => pi,
677 => wh,
678 => wh,
679 => wh,
680 => wh,
681 => wh,
682 => wh,
683 => wh,
684 => sa,
685 => wh,
686 => wh,
687 => wh,
688 => wh,
689 => wh,
690 => wh,
691 => wh,
692 => wh,
693 => wh,
694 => wh,
695 => wh,
696 => wh,
697 => wh,
698 => wh,
699 => pi,
700 => wh,
701 => wh,
702 => wh,
703 => wh,
704 => wh,
705 => wh,
706 => sb,
707 => lb,
708 => lb,
709 => sb,
710 => wh,
711 => wh,
712 => wh,
713 => wh,
714 => pi,
715 => lb,
716 => lb,
717 => sb,
718 => wh,
719 => wh,
720 => wh,
721 => wh,
722 => sb,
723 => lb,
724 => sa,
725 => lb,
726 => sb,
727 => wh,
728 => wh,
729 => wh,
730 => pi,
731 => lb,
732 => sa,
733 => pi,
734 => wh,
735 => wh,
736 => wh,
737 => wh,
738 => sb,
739 => sa,
740 => lb,
741 => sb,
742 => wh,
743 => wh,
744 => wh,
745 => pi,
746 => sa,
747 => lb,
748 => sa,
749 => sb,
750 => wh,
751 => wh,
752 => wh,
753 => wh,
754 => pi,
755 => sa,
756 => sa,
757 => pi,
758 => wh,
759 => wh,
760 => wh,
761 => wh,
762 => pi,
763 => sa,
764 => sa,
765 => pi,
766 => wh,
767 => wh,
768 => wh,
769 => wh,
770 => wh,
771 => wh,
772 => wh,
773 => wh,
774 => wh,
775 => wh,
776 => wh,
777 => wh,
778 => wh,
779 => wh,
780 => wh,
781 => wh,
782 => wh,
783 => wh,
784 => wh,
785 => wh,
786 => wh,
787 => wh,
788 => wh,
789 => wh,
790 => wh,
791 => wh,
792 => wh,
793 => wh,
794 => wh,
795 => wh,
796 => wh,
797 => wh,
798 => wh,
799 => wh,
800 => wh,
801 => wh,
802 => wh,
803 => wh,
804 => wh,
805 => wh,
806 => wh,
807 => dg,
808 => wh,
809 => wh,
810 => wh,
811 => wh,
812 => wh,
813 => wh,
814 => wh,
815 => dg,
816 => wh,
817 => wh,
818 => wh,
819 => wh,
820 => wh,
821 => wh,
822 => dg,
823 => dg,
824 => wh,
825 => wh,
826 => wh,
827 => wh,
828 => wh,
829 => wh,
830 => dg,
831 => ge,
832 => dg,
833 => wh,
834 => wh,
835 => wh,
836 => wh,
837 => wh,
838 => wh,
839 => wh,
840 => dg,
841 => wh,
842 => wh,
843 => wh,
844 => wh,
845 => wh,
846 => wh,
847 => wh,
848 => dg,
849 => wh,
850 => wh,
851 => wh,
852 => wh,
853 => wh,
854 => wh,
855 => wh,
856 => dg,
857 => wh,
858 => wh,
859 => wh,
860 => wh,
861 => wh,
862 => wh,
863 => wh,
864 => wh,
865 => dg,
866 => wh,
867 => wh,
868 => wh,
869 => wh,
870 => wh,
871 => wh,
872 => pi,
873 => pu,
874 => wh,
875 => wh,
876 => wh,
877 => wh,
878 => wh,
879 => wh,
880 => dg,
881 => wh,
882 => dg,
883 => wh,
884 => wh,
885 => wh,
886 => wh,
887 => wh,
888 => dg,
889 => pi,
890 => pu,
891 => wh,
892 => wh,
893 => wh,
894 => wh,
895 => wh,
896 => wh,
897 => wh,
898 => wh,
899 => wh,
900 => wh,
901 => dg,
902 => dg,
903 => wh,
904 => wh,
905 => wh,
906 => wh,
907 => wh,
908 => dg,
909 => dg,
910 => ge,
911 => ge,
912 => wh,
913 => wh,
914 => wh,
915 => wh,
916 => wh,
917 => dg,
918 => dg,
919 => dg,
920 => wh,
921 => wh,
922 => wh,
923 => wh,
924 => dg,
925 => dg,
926 => dg,
927 => wh,
928 => wh,
929 => wh,
930 => wh,
931 => dg,
932 => dg,
933 => dg,
934 => wh,
935 => ge,
936 => wh,
937 => wh,
938 => wh,
939 => wh,
940 => dg,
941 => ge,
942 => ge,
943 => ge,
944 => wh,
945 => wh,
946 => wh,
947 => dg,
948 => dg,
949 => dg,
950 => dg,
951 => pu,
952 => wh,
953 => dg,
954 => dg,
955 => dg,
956 => ge,
957 => wh,
958 => wh,
959 => pi,
960 => ge,
961 => ge,
962 => ge,
963 => pu,
964 => wh,
965 => wh,
966 => wh,
967 => wh,
968 => ge,
969 => ge,
970 => ge,
971 => ge,
972 => dg,
973 => wh,
974 => wh,
975 => wh,
976 => pu,
977 => dg,
978 => pu,
979 => pu,
980 => wh,
981 => wh,
982 => wh,
983 => wh,
984 => pi,
985 => ge,
986 => wh,
987 => pi,
988 => dg,
989 => wh,
990 => wh,
991 => wh,
992 => ge,
993 => ge,
994 => ge,
995 => ge,
996 => ge,
997 => dg,
998 => wh,
999 => wh,
1000 => ge,
1001 => dg,
1002 => pu,
1003 => pu,
1004 => pu,
1005 => wh,
1006 => wh,
1007 => wh,
1008 => dg,
1009 => pu,
1010 => ge,
1011 => wh,
1012 => pi,
1013 => dg,
1014 => wh,
1015 => wh,
1016 => ge,
1017 => pi,
1018 => ge,
1019 => ge,
1020 => ge,
1021 => ge,
1022 => pu,
1023 => dg,
1024 => wh,
1025 => wh,
1026 => pu,
1027 => pu,
1028 => pu,
1029 => pu,
1030 => ge,
1031 => ge,
1032 => wh,
1033 => wh,
1034 => wh,
1035 => pu,
1036 => pu,
1037 => pu,
1038 => pu,
1039 => pu,
1040 => pu,
1041 => pu,
1042 => pu,
1043 => pu,
1044 => ge,
1045 => wh,
1046 => ge,
1047 => wh,
1048 => wh,
1049 => pu,
1050 => pu,
1051 => pu,
1052 => ge,
1053 => ge,
1054 => ge,
1055 => ge,
1056 => wh,
1057 => wh,
1058 => wh,
1059 => wh,
1060 => pu,
1061 => pu,
1062 => ge,
1063 => pu,
1064 => wh,
1065 => wh,
1066 => wh,
1067 => wh,
1068 => wh,
1069 => wh,
1070 => br,
1071 => br,
1072 => wh,
1073 => wh,
1074 => wh,
1075 => wh,
1076 => wh,
1077 => wh,
1078 => lo,
1079 => lo,
1080 => wh,
1081 => wh,
1082 => wh,
1083 => wh,
1084 => wh,
1085 => wh,
1086 => lo,
1087 => lo,
1088 => ge,
1089 => ge,
1090 => ge,
1091 => pu,
1092 => dg,
1093 => pu,
1094 => dg,
1095 => wh,
1096 => pu,
1097 => dg,
1098 => pu,
1099 => pu,
1100 => pu,
1101 => dg,
1102 => wh,
1103 => wh,
1104 => pi,
1105 => pi,
1106 => ge,
1107 => wh,
1108 => pi,
1109 => ge,
1110 => pi,
1111 => pu,
1112 => ge,
1113 => ge,
1114 => ge,
1115 => ge,
1116 => dg,
1117 => dg,
1118 => dg,
1119 => wh,
1120 => dg,
1121 => pu,
1122 => pu,
1123 => dg,
1124 => pu,
1125 => wh,
1126 => wh,
1127 => wh,
1128 => br,
1129 => br,
1130 => br,
1131 => wh,
1132 => wh,
1133 => wh,
1134 => wh,
1135 => wh,
1136 => br,
1137 => br,
1138 => br,
1139 => wh,
1140 => wh,
1141 => wh,
1142 => wh,
1143 => wh,
1144 => lo,
1145 => br,
1146 => br,
1147 => wh,
1148 => wh,
1149 => wh,
1150 => wh,
1151 => wh,
1152 => wh,
1153 => wh,
1154 => wh,
1155 => wh,
1156 => pi,
1157 => wh,
1158 => wh,
1159 => wh,
1160 => wh,
1161 => wh,
1162 => wh,
1163 => ge,
1164 => ge,
1165 => wh,
1166 => wh,
1167 => wh,
1168 => wh,
1169 => wh,
1170 => dg,
1171 => wh,
1172 => ge,
1173 => pi,
1174 => wh,
1175 => wh,
1176 => wh,
1177 => dg,
1178 => ge,
1179 => ge,
1180 => wh,
1181 => dg,
1182 => pu,
1183 => wh,
1184 => wh,
1185 => wh,
1186 => dg,
1187 => dg,
1188 => dg,
1189 => pu,
1190 => wh,
1191 => wh,
1192 => wh,
1193 => pu,
1194 => pu,
1195 => pu,
1196 => pu,
1197 => pu,
1198 => pu,
1199 => wh,
1200 => wh,
1201 => wh,
1202 => wh,
1203 => br,
1204 => br,
1205 => wh,
1206 => wh,
1207 => wh,
1208 => wh,
1209 => wh,
1210 => wh,
1211 => wh,
1212 => wh,
1213 => wh,
1214 => wh,
1215 => wh,
1216 => wh,
1217 => wh,
1218 => wh,
1219 => wh,
1220 => wh,
1221 => wh,
1222 => wh,
1223 => wh,
1224 => wh,
1225 => wh,
1226 => wh,
1227 => ye,
1228 => oa,
1229 => wh,
1230 => wh,
1231 => wh,
1232 => wh,
1233 => wh,
1234 => ye,
1235 => ye,
1236 => ye,
1237 => oa,
1238 => wh,
1239 => wh,
1240 => wh,
1241 => wh,
1242 => ye,
1243 => ye,
1244 => ye,
1245 => oa,
1246 => wh,
1247 => wh,
1248 => wh,
1249 => wh,
1250 => ye,
1251 => ye,
1252 => ye,
1253 => oa,
1254 => wh,
1255 => wh,
1256 => wh,
1257 => wh,
1258 => ye,
1259 => ye,
1260 => ye,
1261 => oa,
1262 => wh,
1263 => wh,
1264 => wh,
1265 => wh,
1266 => wh,
1267 => ye,
1268 => oa,
1269 => wh,
1270 => wh,
1271 => wh,
1272 => wh,
1273 => wh,
1274 => wh,
1275 => wh,
1276 => wh,
1277 => wh,
1278 => wh,
1279 => wh,
1280 => wh,
1281 => wh,
1282 => wh,
1283 => wh,
1284 => wh,
1285 => wh,
1286 => sa,
1287 => wh,
1288 => wh,
1289 => wh,
1290 => wh,
1291 => wh,
1292 => wh,
1293 => sa,
1294 => ye,
1295 => sa,
1296 => wh,
1297 => wh,
1298 => sa,
1299 => wh,
1300 => wh,
1301 => wh,
1302 => sa,
1303 => wh,
1304 => wh,
1305 => sa,
1306 => ye,
1307 => sa,
1308 => wh,
1309 => wh,
1310 => wh,
1311 => wh,
1312 => wh,
1313 => wh,
1314 => sa,
1315 => wh,
1316 => wh,
1317 => sa,
1318 => wh,
1319 => wh,
1320 => wh,
1321 => wh,
1322 => wh,
1323 => wh,
1324 => sa,
1325 => ye,
1326 => sa,
1327 => wh,
1328 => wh,
1329 => wh,
1330 => wh,
1331 => wh,
1332 => wh,
1333 => sa,
1334 => wh,
1335 => wh,
1336 => wh,
1337 => wh,
1338 => wh,
1339 => wh,
1340 => wh,
1341 => wh,
1342 => wh,
1343 => wh,
1344 => wh,
1345 => ye,
1346 => wh,
1347 => wh,
1348 => wh,
1349 => wh,
1350 => wh,
1351 => wh,
1352 => ye,
1353 => oa,
1354 => ye,
1355 => wh,
1356 => wh,
1357 => wh,
1358 => wh,
1359 => wh,
1360 => wh,
1361 => ye,
1362 => wh,
1363 => wh,
1364 => wh,
1365 => ye,
1366 => wh,
1367 => wh,
1368 => wh,
1369 => wh,
1370 => wh,
1371 => wh,
1372 => ye,
1373 => oa,
1374 => ye,
1375 => wh,
1376 => wh,
1377 => wh,
1378 => ye,
1379 => wh,
1380 => wh,
1381 => ye,
1382 => wh,
1383 => wh,
1384 => wh,
1385 => ye,
1386 => oa,
1387 => ye,
1388 => wh,
1389 => wh,
1390 => wh,
1391 => wh,
1392 => wh,
1393 => wh,
1394 => ye,
1395 => wh,
1396 => wh,
1397 => wh,
1398 => wh,
1399 => wh,
1400 => wh,
1401 => wh,
1402 => wh,
1403 => wh,
1404 => wh,
1405 => wh,
1406 => wh,
1407 => wh,
1408 => wh,
1409 => pi,
1410 => lg,
1411 => wh,
1412 => wh,
1413 => wh,
1414 => wh,
1415 => wh,
1416 => wh,
1417 => lg,
1418 => lg,
1419 => lo,
1420 => lo,
1421 => lo,
1422 => lo,
1423 => br,
1424 => wh,
1425 => lg,
1426 => gr,
1427 => br,
1428 => br,
1429 => br,
1430 => br,
1431 => br,
1432 => wh,
1433 => lg,
1434 => lg,
1435 => wh,
1436 => wh,
1437 => wh,
1438 => wh,
1439 => wh,
1440 => wh,
1441 => gr,
1442 => gr,
1443 => lo,
1444 => lo,
1445 => br,
1446 => br,
1447 => lo,
1448 => wh,
1449 => lg,
1450 => gr,
1451 => lo,
1452 => lo,
1453 => lo,
1454 => lo,
1455 => lo,
1456 => wh,
1457 => gr,
1458 => lg,
1459 => br,
1460 => br,
1461 => br,
1462 => br,
1463 => pi,
1464 => wh,
1465 => gr,
1466 => pi,
1467 => wh,
1468 => wh,
1469 => wh,
1470 => wh,
1471 => wh,
1472 => wh,
1473 => wh,
1474 => wh,
1475 => wh,
1476 => wh,
1477 => wh,
1478 => wh,
1479 => wh,
1480 => lo,
1481 => lo,
1482 => lo,
1483 => lo,
1484 => lo,
1485 => br,
1486 => lo,
1487 => lo,
1488 => br,
1489 => br,
1490 => br,
1491 => br,
1492 => br,
1493 => pi,
1494 => br,
1495 => br,
1496 => wh,
1497 => wh,
1498 => wh,
1499 => wh,
1500 => wh,
1501 => wh,
1502 => wh,
1503 => wh,
1504 => lo,
1505 => lo,
1506 => lo,
1507 => pi,
1508 => lo,
1509 => lo,
1510 => lo,
1511 => lo,
1512 => br,
1513 => lo,
1514 => lo,
1515 => br,
1516 => lo,
1517 => br,
1518 => lo,
1519 => lo,
1520 => br,
1521 => wh,
1522 => wh,
1523 => br,
1524 => br,
1525 => br,
1526 => br,
1527 => br,
1528 => wh,
1529 => wh,
1530 => wh,
1531 => wh,
1532 => wh,
1533 => wh,
1534 => wh,
1535 => wh,
        others => bl
    ); 
    
    attribute ram_style : string;
    attribute ram_style of tile_data_map_d : signal is "block";
begin
    
      process(i_tile_id, i_x, i_y)
          variable readIndex : std_logic_vector (10 downto 0);
          variable readIndex_int : integer;
          begin
          readIndex := i_tile_id & i_y & i_x;
          readIndex_int := to_integer(unsigned(readIndex));
          o_colorCode <= tile_data_map_d(readIndex_int);
      end process;
      
      process(i_clk)
      variable writeIndex : std_logic_vector (10 downto 0);
      variable writeIndex_int : integer;
      begin
        if rising_edge(i_clk) then
            if i_ch_we = '1' then
                writeIndex := i_tile_id_write & i_ch_y & i_ch_x;
                writeIndex_int := to_integer(unsigned(writeIndex));
                tile_data_map_d(writeIndex_int) <= i_ch_cc;
            end if;
        end if;
      end process;

end Behavioral;
