----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08.06.2025 00:00:57
-- Design Name: 
-- Module Name: BackMgmt - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity BackMgmt is
    Port ( 
        i_view_x : in STD_LOGIC_VECTOR (9 downto 0); -- position x du pixel � voir
        i_view_y : in STD_LOGIC_VECTOR (9 downto 0); -- position y du pixel � voir
        i_ch_we_tileBack : in STD_LOGIC;
        i_col : in STD_LOGIC_VECTOR (6 downto 0); -- prochaine tuile � changer
        i_row : in STD_LOGIC_VECTOR (6 downto 0); -- prochaine tuile � changer
        i_tile_id : in STD_LOGIC_VECTOR (4 downto 0); -- tuile qui change
        i_flip_y : in STD_LOGIC; -- valeur du flip
        i_ch_tile_id : in STD_LOGIC; -- change la tuile?
        i_ch_flip_y : in STD_LOGIC; -- change le flip?
        i_clk : in STD_LOGIC; -- la clock

        -- Info du pixel qu'on regarde
        o_tile_id : out STD_LOGIC_VECTOR (4 downto 0); 
        o_flip_y : out STD_LOGIC;
        o_pix_x : out STD_LOGIC_VECTOR (2 downto 0);
        o_pix_y : out STD_LOGIC_VECTOR (2 downto 0)
    );
end BackMgmt;

architecture Behavioral of BackMgmt is

    -- Packed format: [5] = flip_y, [4:0] = tile_id
    type tile_data_array_t is array (0 to 16383) of std_logic_vector(7 downto 0);
    signal tile_data_map : tile_data_array_t := (
        1 => "00000010",
129 => "00000010",
257 => "00000010",
385 => "00000010",
513 => "00000010",
641 => "00000010",
769 => "00000010",
897 => "00000010",
1025 => "00000010",
1153 => "00000010",
1281 => "00000010",
1409 => "00000010",
1537 => "00000010",
1665 => "00000010",
1793 => "00000010",
1921 => "00000010",
2049 => "00000010",
2177 => "00000010",
2305 => "00000010",
2433 => "00000010",
2561 => "00000010",
2689 => "00000010",
2817 => "00000010",
2945 => "00000010",
3073 => "00000010",
3201 => "00000010",
3329 => "00000010",
3457 => "00000010",
3585 => "00000010",
3713 => "00000010",
3841 => "00000010",
3969 => "00000010",
4097 => "00000010",
4225 => "00000010",
4353 => "00000010",
4481 => "00000010",
4609 => "00000010",
4737 => "00000010",
4865 => "00000010",
4993 => "00000010",
5121 => "00000010",
5249 => "00000010",
5377 => "00000010",
5505 => "00000010",
5633 => "00000010",
5761 => "00000010",
5889 => "00000010",
6017 => "00000010",
6145 => "00000010",
6273 => "00000010",
6401 => "00000010",
6529 => "00000010",
6657 => "00000010",
6785 => "00000010",
6913 => "00000010",
7041 => "00000010",
7169 => "00000010",
7297 => "00000010",
7425 => "00000010",
7553 => "00000010",
7681 => "00000010",
7809 => "00000010",
7937 => "00000010",
8065 => "00000010",
8193 => "00000010",
8321 => "00000010",
8449 => "00000010",
8577 => "00000010",
8705 => "00000010",
8833 => "00000010",
8961 => "00000010",
9089 => "00000010",
9217 => "00000010",
9345 => "00000010",
9473 => "00000010",
9601 => "00000010",
9729 => "00000010",
9857 => "00000010",
9985 => "00000010",
10113 => "00000010",
10241 => "00000010",
10369 => "00000010",
10497 => "00000010",
10625 => "00000010",
10753 => "00000010",
10881 => "00000010",
11009 => "00000010",
11137 => "00000010",
11265 => "00000010",
11393 => "00000010",
11521 => "00000010",
11649 => "00000010",
11777 => "00000010",
11905 => "00000010",
12033 => "00000010",
12161 => "00000010",
12289 => "00000010",
12417 => "00000010",
12545 => "00000010",
12673 => "00000010",
12801 => "00000010",
12929 => "00000010",
13057 => "00000010",
13185 => "00000010",
13313 => "00000010",
13441 => "00000010",
13569 => "00000010",
13697 => "00000010",
13825 => "00000010",
13953 => "00000010",
14081 => "00000010",
14209 => "00000010",
14337 => "00000010",
14465 => "00000010",
14593 => "00000010",
14721 => "00000010",
14849 => "00000010",
14977 => "00000010",
15105 => "00000010",
15233 => "00000010",
15361 => "00000010",
15489 => "00000010",
15617 => "00000010",
15745 => "00000010",
15873 => "00000010",
16001 => "00000010",
16129 => "00000010",
16257 => "00000010",
7 => "00000001",
135 => "00000001",
263 => "00000001",
391 => "00000001",
519 => "00000001",
647 => "00000001",
775 => "00000001",
903 => "00000001",
1031 => "00000001",
1159 => "00000001",
1287 => "00000001",
1415 => "00000001",
1543 => "00000001",
1671 => "00000001",
1799 => "00000001",
1927 => "00000001",
2055 => "00000001",
2183 => "00000001",
2311 => "00000001",
2439 => "00000001",
2567 => "00000001",
2695 => "00000001",
2823 => "00000001",
2951 => "00000001",
3079 => "00000001",
3207 => "00000001",
3335 => "00000001",
3463 => "00000001",
3591 => "00000001",
3719 => "00000001",
3847 => "00000001",
3975 => "00000001",
4103 => "00000001",
4231 => "00000001",
4359 => "00000001",
4487 => "00000001",
4615 => "00000001",
4743 => "00000001",
4871 => "00000001",
4999 => "00000001",
5127 => "00000001",
5255 => "00000001",
5383 => "00000001",
5511 => "00000001",
5639 => "00000001",
5767 => "00000001",
5895 => "00000001",
6023 => "00000001",
6151 => "00000001",
6279 => "00000001",
6407 => "00000001",
6535 => "00000001",
6663 => "00000001",
6791 => "00000001",
6919 => "00000001",
7047 => "00000001",
7175 => "00000001",
7303 => "00000001",
7431 => "00000001",
7559 => "00000001",
7687 => "00000001",
7815 => "00000001",
7943 => "00000001",
8071 => "00000001",
8199 => "00000001",
8327 => "00000001",
8455 => "00000001",
8583 => "00000001",
8711 => "00000001",
8839 => "00000001",
8967 => "00000001",
9095 => "00000001",
9223 => "00000001",
9351 => "00000001",
9479 => "00000001",
9607 => "00000001",
9735 => "00000001",
9863 => "00000001",
9991 => "00000001",
10119 => "00000001",
10247 => "00000001",
10375 => "00000001",
10503 => "00000001",
10631 => "00000001",
10759 => "00000001",
10887 => "00000001",
11015 => "00000001",
11143 => "00000001",
11271 => "00000001",
11399 => "00000001",
11527 => "00000001",
11655 => "00000001",
11783 => "00000001",
11911 => "00000001",
12039 => "00000001",
12167 => "00000001",
12295 => "00000001",
12423 => "00000001",
12551 => "00000001",
12679 => "00000001",
12807 => "00000001",
12935 => "00000001",
13063 => "00000001",
13191 => "00000001",
13319 => "00000001",
13447 => "00000001",
13575 => "00000001",
13703 => "00000001",
13831 => "00000001",
13959 => "00000001",
14087 => "00000001",
14215 => "00000001",
14343 => "00000001",
14471 => "00000001",
14599 => "00000001",
14727 => "00000001",
14855 => "00000001",
14983 => "00000001",
15111 => "00000001",
15239 => "00000001",
15367 => "00000001",
15495 => "00000001",
15623 => "00000001",
15751 => "00000001",
15879 => "00000001",
16007 => "00000001",
16135 => "00000001",
16263 => "00000001",
13 => "00000001",
141 => "00000001",
269 => "00000001",
397 => "00000001",
525 => "00000001",
653 => "00000001",
781 => "00000001",
909 => "00000001",
1037 => "00000001",
1165 => "00000001",
1293 => "00000001",
1421 => "00000001",
1549 => "00000001",
1677 => "00000001",
1805 => "00000001",
1933 => "00000001",
2061 => "00000001",
2189 => "00000001",
2317 => "00000001",
2445 => "00000001",
2573 => "00000001",
2701 => "00000001",
2829 => "00000001",
2957 => "00000001",
3085 => "00000001",
3213 => "00000001",
3341 => "00000001",
3469 => "00000001",
3597 => "00000001",
3725 => "00000001",
3853 => "00000001",
3981 => "00000001",
4109 => "00000001",
4237 => "00000001",
4365 => "00000001",
4493 => "00000001",
4621 => "00000001",
4749 => "00000001",
4877 => "00000001",
5005 => "00000001",
5133 => "00000001",
5261 => "00000001",
5389 => "00000001",
5517 => "00000001",
5645 => "00000001",
5773 => "00000001",
5901 => "00000001",
6029 => "00000001",
6157 => "00000001",
6285 => "00000001",
6413 => "00000001",
6541 => "00000001",
6669 => "00000001",
6797 => "00000001",
6925 => "00000001",
7053 => "00000001",
7181 => "00000001",
7309 => "00000001",
7437 => "00000001",
7565 => "00000001",
7693 => "00000001",
7821 => "00000001",
7949 => "00000001",
8077 => "00000001",
8205 => "00000001",
8333 => "00000001",
8461 => "00000001",
8589 => "00000001",
8717 => "00000001",
8845 => "00000001",
8973 => "00000001",
9101 => "00000001",
9229 => "00000001",
9357 => "00000001",
9485 => "00000001",
9613 => "00000001",
9741 => "00000001",
9869 => "00000001",
9997 => "00000001",
10125 => "00000001",
10253 => "00000001",
10381 => "00000001",
10509 => "00000001",
10637 => "00000001",
10765 => "00000001",
10893 => "00000001",
11021 => "00000001",
11149 => "00000001",
11277 => "00000001",
11405 => "00000001",
11533 => "00000001",
11661 => "00000001",
11789 => "00000001",
11917 => "00000001",
12045 => "00000001",
12173 => "00000001",
12301 => "00000001",
12429 => "00000001",
12557 => "00000001",
12685 => "00000001",
12813 => "00000001",
12941 => "00000001",
13069 => "00000001",
13197 => "00000001",
13325 => "00000001",
13453 => "00000001",
13581 => "00000001",
13709 => "00000001",
13837 => "00000001",
13965 => "00000001",
14093 => "00000001",
14221 => "00000001",
14349 => "00000001",
14477 => "00000001",
14605 => "00000001",
14733 => "00000001",
14861 => "00000001",
14989 => "00000001",
15117 => "00000001",
15245 => "00000001",
15373 => "00000001",
15501 => "00000001",
15629 => "00000001",
15757 => "00000001",
15885 => "00000001",
16013 => "00000001",
16141 => "00000001",
16269 => "00000001",
19 => "00000001",
147 => "00000001",
275 => "00000001",
403 => "00000001",
531 => "00000001",
659 => "00000001",
787 => "00000001",
915 => "00000001",
1043 => "00000001",
1171 => "00000001",
1299 => "00000001",
1427 => "00000001",
1555 => "00000001",
1683 => "00000001",
1811 => "00000001",
1939 => "00000001",
2067 => "00000001",
2195 => "00000001",
2323 => "00000001",
2451 => "00000001",
2579 => "00000001",
2707 => "00000001",
2835 => "00000001",
2963 => "00000001",
3091 => "00000001",
3219 => "00000001",
3347 => "00000001",
3475 => "00000001",
3603 => "00000001",
3731 => "00000001",
3859 => "00000001",
3987 => "00000001",
4115 => "00000001",
4243 => "00000001",
4371 => "00000001",
4499 => "00000001",
4627 => "00000001",
4755 => "00000001",
4883 => "00000001",
5011 => "00000001",
5139 => "00000001",
5267 => "00000001",
5395 => "00000001",
5523 => "00000001",
5651 => "00000001",
5779 => "00000001",
5907 => "00000001",
6035 => "00000001",
6163 => "00000001",
6291 => "00000001",
6419 => "00000001",
6547 => "00000001",
6675 => "00000001",
6803 => "00000001",
6931 => "00000001",
7059 => "00000001",
7187 => "00000001",
7315 => "00000001",
7443 => "00000001",
7571 => "00000001",
7699 => "00000001",
7827 => "00000001",
7955 => "00000001",
8083 => "00000001",
8211 => "00000001",
8339 => "00000001",
8467 => "00000001",
8595 => "00000001",
8723 => "00000001",
8851 => "00000001",
8979 => "00000001",
9107 => "00000001",
9235 => "00000001",
9363 => "00000001",
9491 => "00000001",
9619 => "00000001",
9747 => "00000001",
9875 => "00000001",
10003 => "00000001",
10131 => "00000001",
10259 => "00000001",
10387 => "00000001",
10515 => "00000001",
10643 => "00000001",
10771 => "00000001",
10899 => "00000001",
11027 => "00000001",
11155 => "00000001",
11283 => "00000001",
11411 => "00000001",
11539 => "00000001",
11667 => "00000001",
11795 => "00000001",
11923 => "00000001",
12051 => "00000001",
12179 => "00000001",
12307 => "00000001",
12435 => "00000001",
12563 => "00000001",
12691 => "00000001",
12819 => "00000001",
12947 => "00000001",
13075 => "00000001",
13203 => "00000001",
13331 => "00000001",
13459 => "00000001",
13587 => "00000001",
13715 => "00000001",
13843 => "00000001",
13971 => "00000001",
14099 => "00000001",
14227 => "00000001",
14355 => "00000001",
14483 => "00000001",
14611 => "00000001",
14739 => "00000001",
14867 => "00000001",
14995 => "00000001",
15123 => "00000001",
15251 => "00000001",
15379 => "00000001",
15507 => "00000001",
15635 => "00000001",
15763 => "00000001",
15891 => "00000001",
16019 => "00000001",
16147 => "00000001",
16275 => "00000001",
25 => "00000001",
153 => "00000001",
281 => "00000001",
409 => "00000001",
537 => "00000001",
665 => "00000001",
793 => "00000001",
921 => "00000001",
1049 => "00000001",
1177 => "00000001",
1305 => "00000001",
1433 => "00000001",
1561 => "00000001",
1689 => "00000001",
1817 => "00000001",
1945 => "00000001",
2073 => "00000001",
2201 => "00000001",
2329 => "00000001",
2457 => "00000001",
2585 => "00000001",
2713 => "00000001",
2841 => "00000001",
2969 => "00000001",
3097 => "00000001",
3225 => "00000001",
3353 => "00000001",
3481 => "00000001",
3609 => "00000001",
3737 => "00000001",
3865 => "00000001",
3993 => "00000001",
4121 => "00000001",
4249 => "00000001",
4377 => "00000001",
4505 => "00000001",
4633 => "00000001",
4761 => "00000001",
4889 => "00000001",
5017 => "00000001",
5145 => "00000001",
5273 => "00000001",
5401 => "00000001",
5529 => "00000001",
5657 => "00000001",
5785 => "00000001",
5913 => "00000001",
6041 => "00000001",
6169 => "00000001",
6297 => "00000001",
6425 => "00000001",
6553 => "00000001",
6681 => "00000001",
6809 => "00000001",
6937 => "00000001",
7065 => "00000001",
7193 => "00000001",
7321 => "00000001",
7449 => "00000001",
7577 => "00000001",
7705 => "00000001",
7833 => "00000001",
7961 => "00000001",
8089 => "00000001",
8217 => "00000001",
8345 => "00000001",
8473 => "00000001",
8601 => "00000001",
8729 => "00000001",
8857 => "00000001",
8985 => "00000001",
9113 => "00000001",
9241 => "00000001",
9369 => "00000001",
9497 => "00000001",
9625 => "00000001",
9753 => "00000001",
9881 => "00000001",
10009 => "00000001",
10137 => "00000001",
10265 => "00000001",
10393 => "00000001",
10521 => "00000001",
10649 => "00000001",
10777 => "00000001",
10905 => "00000001",
11033 => "00000001",
11161 => "00000001",
11289 => "00000001",
11417 => "00000001",
11545 => "00000001",
11673 => "00000001",
11801 => "00000001",
11929 => "00000001",
12057 => "00000001",
12185 => "00000001",
12313 => "00000001",
12441 => "00000001",
12569 => "00000001",
12697 => "00000001",
12825 => "00000001",
12953 => "00000001",
13081 => "00000001",
13209 => "00000001",
13337 => "00000001",
13465 => "00000001",
13593 => "00000001",
13721 => "00000001",
13849 => "00000001",
13977 => "00000001",
14105 => "00000001",
14233 => "00000001",
14361 => "00000001",
14489 => "00000001",
14617 => "00000001",
14745 => "00000001",
14873 => "00000001",
15001 => "00000001",
15129 => "00000001",
15257 => "00000001",
15385 => "00000001",
15513 => "00000001",
15641 => "00000001",
15769 => "00000001",
15897 => "00000001",
16025 => "00000001",
16153 => "00000001",
16281 => "00000001",
31 => "00000001",
159 => "00000001",
287 => "00000001",
415 => "00000001",
543 => "00000001",
671 => "00000001",
799 => "00000001",
927 => "00000001",
1055 => "00000001",
1183 => "00000001",
1311 => "00000001",
1439 => "00000001",
1567 => "00000001",
1695 => "00000001",
1823 => "00000001",
1951 => "00000001",
2079 => "00000001",
2207 => "00000001",
2335 => "00000001",
2463 => "00000001",
2591 => "00000001",
2719 => "00000001",
2847 => "00000001",
2975 => "00000001",
3103 => "00000001",
3231 => "00000001",
3359 => "00000001",
3487 => "00000001",
3615 => "00000001",
3743 => "00000001",
3871 => "00000001",
3999 => "00000001",
4127 => "00000001",
4255 => "00000001",
4383 => "00000001",
4511 => "00000001",
4639 => "00000001",
4767 => "00000001",
4895 => "00000001",
5023 => "00000001",
5151 => "00000001",
5279 => "00000001",
5407 => "00000001",
5535 => "00000001",
5663 => "00000001",
5791 => "00000001",
5919 => "00000001",
6047 => "00000001",
6175 => "00000001",
6303 => "00000001",
6431 => "00000001",
6559 => "00000001",
6687 => "00000001",
6815 => "00000001",
6943 => "00000001",
7071 => "00000001",
7199 => "00000001",
7327 => "00000001",
7455 => "00000001",
7583 => "00000001",
7711 => "00000001",
7839 => "00000001",
7967 => "00000001",
8095 => "00000001",
8223 => "00000001",
8351 => "00000001",
8479 => "00000001",
8607 => "00000001",
8735 => "00000001",
8863 => "00000001",
8991 => "00000001",
9119 => "00000001",
9247 => "00000001",
9375 => "00000001",
9503 => "00000001",
9631 => "00000001",
9759 => "00000001",
9887 => "00000001",
10015 => "00000001",
10143 => "00000001",
10271 => "00000001",
10399 => "00000001",
10527 => "00000001",
10655 => "00000001",
10783 => "00000001",
10911 => "00000001",
11039 => "00000001",
11167 => "00000001",
11295 => "00000001",
11423 => "00000001",
11551 => "00000001",
11679 => "00000001",
11807 => "00000001",
11935 => "00000001",
12063 => "00000001",
12191 => "00000001",
12319 => "00000001",
12447 => "00000001",
12575 => "00000001",
12703 => "00000001",
12831 => "00000001",
12959 => "00000001",
13087 => "00000001",
13215 => "00000001",
13343 => "00000001",
13471 => "00000001",
13599 => "00000001",
13727 => "00000001",
13855 => "00000001",
13983 => "00000001",
14111 => "00000001",
14239 => "00000001",
14367 => "00000001",
14495 => "00000001",
14623 => "00000001",
14751 => "00000001",
14879 => "00000001",
15007 => "00000001",
15135 => "00000001",
15263 => "00000001",
15391 => "00000001",
15519 => "00000001",
15647 => "00000001",
15775 => "00000001",
15903 => "00000001",
16031 => "00000001",
16159 => "00000001",
16287 => "00000001",
37 => "00000001",
165 => "00000001",
293 => "00000001",
421 => "00000001",
549 => "00000001",
677 => "00000001",
805 => "00000001",
933 => "00000001",
1061 => "00000001",
1189 => "00000001",
1317 => "00000001",
1445 => "00000001",
1573 => "00000001",
1701 => "00000001",
1829 => "00000001",
1957 => "00000001",
2085 => "00000001",
2213 => "00000001",
2341 => "00000001",
2469 => "00000001",
2597 => "00000001",
2725 => "00000001",
2853 => "00000001",
2981 => "00000001",
3109 => "00000001",
3237 => "00000001",
3365 => "00000001",
3493 => "00000001",
3621 => "00000001",
3749 => "00000001",
3877 => "00000001",
4005 => "00000001",
4133 => "00000001",
4261 => "00000001",
4389 => "00000001",
4517 => "00000001",
4645 => "00000001",
4773 => "00000001",
4901 => "00000001",
5029 => "00000001",
5157 => "00000001",
5285 => "00000001",
5413 => "00000001",
5541 => "00000001",
5669 => "00000001",
5797 => "00000001",
5925 => "00000001",
6053 => "00000001",
6181 => "00000001",
6309 => "00000001",
6437 => "00000001",
6565 => "00000001",
6693 => "00000001",
6821 => "00000001",
6949 => "00000001",
7077 => "00000001",
7205 => "00000001",
7333 => "00000001",
7461 => "00000001",
7589 => "00000001",
7717 => "00000001",
7845 => "00000001",
7973 => "00000001",
8101 => "00000001",
8229 => "00000001",
8357 => "00000001",
8485 => "00000001",
8613 => "00000001",
8741 => "00000001",
8869 => "00000001",
8997 => "00000001",
9125 => "00000001",
9253 => "00000001",
9381 => "00000001",
9509 => "00000001",
9637 => "00000001",
9765 => "00000001",
9893 => "00000001",
10021 => "00000001",
10149 => "00000001",
10277 => "00000001",
10405 => "00000001",
10533 => "00000001",
10661 => "00000001",
10789 => "00000001",
10917 => "00000001",
11045 => "00000001",
11173 => "00000001",
11301 => "00000001",
11429 => "00000001",
11557 => "00000001",
11685 => "00000001",
11813 => "00000001",
11941 => "00000001",
12069 => "00000001",
12197 => "00000001",
12325 => "00000001",
12453 => "00000001",
12581 => "00000001",
12709 => "00000001",
12837 => "00000001",
12965 => "00000001",
13093 => "00000001",
13221 => "00000001",
13349 => "00000001",
13477 => "00000001",
13605 => "00000001",
13733 => "00000001",
13861 => "00000001",
13989 => "00000001",
14117 => "00000001",
14245 => "00000001",
14373 => "00000001",
14501 => "00000001",
14629 => "00000001",
14757 => "00000001",
14885 => "00000001",
15013 => "00000001",
15141 => "00000001",
15269 => "00000001",
15397 => "00000001",
15525 => "00000001",
15653 => "00000001",
15781 => "00000001",
15909 => "00000001",
16037 => "00000001",
16165 => "00000001",
16293 => "00000001",
43 => "00000001",
171 => "00000001",
299 => "00000001",
427 => "00000001",
555 => "00000001",
683 => "00000001",
811 => "00000001",
939 => "00000001",
1067 => "00000001",
1195 => "00000001",
1323 => "00000001",
1451 => "00000001",
1579 => "00000001",
1707 => "00000001",
1835 => "00000001",
1963 => "00000001",
2091 => "00000001",
2219 => "00000001",
2347 => "00000001",
2475 => "00000001",
2603 => "00000001",
2731 => "00000001",
2859 => "00000001",
2987 => "00000001",
3115 => "00000001",
3243 => "00000001",
3371 => "00000001",
3499 => "00000001",
3627 => "00000001",
3755 => "00000001",
3883 => "00000001",
4011 => "00000001",
4139 => "00000001",
4267 => "00000001",
4395 => "00000001",
4523 => "00000001",
4651 => "00000001",
4779 => "00000001",
4907 => "00000001",
5035 => "00000001",
5163 => "00000001",
5291 => "00000001",
5419 => "00000001",
5547 => "00000001",
5675 => "00000001",
5803 => "00000001",
5931 => "00000001",
6059 => "00000001",
6187 => "00000001",
6315 => "00000001",
6443 => "00000001",
6571 => "00000001",
6699 => "00000001",
6827 => "00000001",
6955 => "00000001",
7083 => "00000001",
7211 => "00000001",
7339 => "00000001",
7467 => "00000001",
7595 => "00000001",
7723 => "00000001",
7851 => "00000001",
7979 => "00000001",
8107 => "00000001",
8235 => "00000001",
8363 => "00000001",
8491 => "00000001",
8619 => "00000001",
8747 => "00000001",
8875 => "00000001",
9003 => "00000001",
9131 => "00000001",
9259 => "00000001",
9387 => "00000001",
9515 => "00000001",
9643 => "00000001",
9771 => "00000001",
9899 => "00000001",
10027 => "00000001",
10155 => "00000001",
10283 => "00000001",
10411 => "00000001",
10539 => "00000001",
10667 => "00000001",
10795 => "00000001",
10923 => "00000001",
11051 => "00000001",
11179 => "00000001",
11307 => "00000001",
11435 => "00000001",
11563 => "00000001",
11691 => "00000001",
11819 => "00000001",
11947 => "00000001",
12075 => "00000001",
12203 => "00000001",
12331 => "00000001",
12459 => "00000001",
12587 => "00000001",
12715 => "00000001",
12843 => "00000001",
12971 => "00000001",
13099 => "00000001",
13227 => "00000001",
13355 => "00000001",
13483 => "00000001",
13611 => "00000001",
13739 => "00000001",
13867 => "00000001",
13995 => "00000001",
14123 => "00000001",
14251 => "00000001",
14379 => "00000001",
14507 => "00000001",
14635 => "00000001",
14763 => "00000001",
14891 => "00000001",
15019 => "00000001",
15147 => "00000001",
15275 => "00000001",
15403 => "00000001",
15531 => "00000001",
15659 => "00000001",
15787 => "00000001",
15915 => "00000001",
16043 => "00000001",
16171 => "00000001",
16299 => "00000001",
49 => "00000001",
177 => "00000001",
305 => "00000001",
433 => "00000001",
561 => "00000001",
689 => "00000001",
817 => "00000001",
945 => "00000001",
1073 => "00000001",
1201 => "00000001",
1329 => "00000001",
1457 => "00000001",
1585 => "00000001",
1713 => "00000001",
1841 => "00000001",
1969 => "00000001",
2097 => "00000001",
2225 => "00000001",
2353 => "00000001",
2481 => "00000001",
2609 => "00000001",
2737 => "00000001",
2865 => "00000001",
2993 => "00000001",
3121 => "00000001",
3249 => "00000001",
3377 => "00000001",
3505 => "00000001",
3633 => "00000001",
3761 => "00000001",
3889 => "00000001",
4017 => "00000001",
4145 => "00000001",
4273 => "00000001",
4401 => "00000001",
4529 => "00000001",
4657 => "00000001",
4785 => "00000001",
4913 => "00000001",
5041 => "00000001",
5169 => "00000001",
5297 => "00000001",
5425 => "00000001",
5553 => "00000001",
5681 => "00000001",
5809 => "00000001",
5937 => "00000001",
6065 => "00000001",
6193 => "00000001",
6321 => "00000001",
6449 => "00000001",
6577 => "00000001",
6705 => "00000001",
6833 => "00000001",
6961 => "00000001",
7089 => "00000001",
7217 => "00000001",
7345 => "00000001",
7473 => "00000001",
7601 => "00000001",
7729 => "00000001",
7857 => "00000001",
7985 => "00000001",
8113 => "00000001",
8241 => "00000001",
8369 => "00000001",
8497 => "00000001",
8625 => "00000001",
8753 => "00000001",
8881 => "00000001",
9009 => "00000001",
9137 => "00000001",
9265 => "00000001",
9393 => "00000001",
9521 => "00000001",
9649 => "00000001",
9777 => "00000001",
9905 => "00000001",
10033 => "00000001",
10161 => "00000001",
10289 => "00000001",
10417 => "00000001",
10545 => "00000001",
10673 => "00000001",
10801 => "00000001",
10929 => "00000001",
11057 => "00000001",
11185 => "00000001",
11313 => "00000001",
11441 => "00000001",
11569 => "00000001",
11697 => "00000001",
11825 => "00000001",
11953 => "00000001",
12081 => "00000001",
12209 => "00000001",
12337 => "00000001",
12465 => "00000001",
12593 => "00000001",
12721 => "00000001",
12849 => "00000001",
12977 => "00000001",
13105 => "00000001",
13233 => "00000001",
13361 => "00000001",
13489 => "00000001",
13617 => "00000001",
13745 => "00000001",
13873 => "00000001",
14001 => "00000001",
14129 => "00000001",
14257 => "00000001",
14385 => "00000001",
14513 => "00000001",
14641 => "00000001",
14769 => "00000001",
14897 => "00000001",
15025 => "00000001",
15153 => "00000001",
15281 => "00000001",
15409 => "00000001",
15537 => "00000001",
15665 => "00000001",
15793 => "00000001",
15921 => "00000001",
16049 => "00000001",
16177 => "00000001",
16305 => "00000001",
55 => "00000001",
183 => "00000001",
311 => "00000001",
439 => "00000001",
567 => "00000001",
695 => "00000001",
823 => "00000001",
951 => "00000001",
1079 => "00000001",
1207 => "00000001",
1335 => "00000001",
1463 => "00000001",
1591 => "00000001",
1719 => "00000001",
1847 => "00000001",
1975 => "00000001",
2103 => "00000001",
2231 => "00000001",
2359 => "00000001",
2487 => "00000001",
2615 => "00000001",
2743 => "00000001",
2871 => "00000001",
2999 => "00000001",
3127 => "00000001",
3255 => "00000001",
3383 => "00000001",
3511 => "00000001",
3639 => "00000001",
3767 => "00000001",
3895 => "00000001",
4023 => "00000001",
4151 => "00000001",
4279 => "00000001",
4407 => "00000001",
4535 => "00000001",
4663 => "00000001",
4791 => "00000001",
4919 => "00000001",
5047 => "00000001",
5175 => "00000001",
5303 => "00000001",
5431 => "00000001",
5559 => "00000001",
5687 => "00000001",
5815 => "00000001",
5943 => "00000001",
6071 => "00000001",
6199 => "00000001",
6327 => "00000001",
6455 => "00000001",
6583 => "00000001",
6711 => "00000001",
6839 => "00000001",
6967 => "00000001",
7095 => "00000001",
7223 => "00000001",
7351 => "00000001",
7479 => "00000001",
7607 => "00000001",
7735 => "00000001",
7863 => "00000001",
7991 => "00000001",
8119 => "00000001",
8247 => "00000001",
8375 => "00000001",
8503 => "00000001",
8631 => "00000001",
8759 => "00000001",
8887 => "00000001",
9015 => "00000001",
9143 => "00000001",
9271 => "00000001",
9399 => "00000001",
9527 => "00000001",
9655 => "00000001",
9783 => "00000001",
9911 => "00000001",
10039 => "00000001",
10167 => "00000001",
10295 => "00000001",
10423 => "00000001",
10551 => "00000001",
10679 => "00000001",
10807 => "00000001",
10935 => "00000001",
11063 => "00000001",
11191 => "00000001",
11319 => "00000001",
11447 => "00000001",
11575 => "00000001",
11703 => "00000001",
11831 => "00000001",
11959 => "00000001",
12087 => "00000001",
12215 => "00000001",
12343 => "00000001",
12471 => "00000001",
12599 => "00000001",
12727 => "00000001",
12855 => "00000001",
12983 => "00000001",
13111 => "00000001",
13239 => "00000001",
13367 => "00000001",
13495 => "00000001",
13623 => "00000001",
13751 => "00000001",
13879 => "00000001",
14007 => "00000001",
14135 => "00000001",
14263 => "00000001",
14391 => "00000001",
14519 => "00000001",
14647 => "00000001",
14775 => "00000001",
14903 => "00000001",
15031 => "00000001",
15159 => "00000001",
15287 => "00000001",
15415 => "00000001",
15543 => "00000001",
15671 => "00000001",
15799 => "00000001",
15927 => "00000001",
16055 => "00000001",
16183 => "00000001",
16311 => "00000001",
61 => "00000001",
189 => "00000001",
317 => "00000001",
445 => "00000001",
573 => "00000001",
701 => "00000001",
829 => "00000001",
957 => "00000001",
1085 => "00000001",
1213 => "00000001",
1341 => "00000001",
1469 => "00000001",
1597 => "00000001",
1725 => "00000001",
1853 => "00000001",
1981 => "00000001",
2109 => "00000001",
2237 => "00000001",
2365 => "00000001",
2493 => "00000001",
2621 => "00000001",
2749 => "00000001",
2877 => "00000001",
3005 => "00000001",
3133 => "00000001",
3261 => "00000001",
3389 => "00000001",
3517 => "00000001",
3645 => "00000001",
3773 => "00000001",
3901 => "00000001",
4029 => "00000001",
4157 => "00000001",
4285 => "00000001",
4413 => "00000001",
4541 => "00000001",
4669 => "00000001",
4797 => "00000001",
4925 => "00000001",
5053 => "00000001",
5181 => "00000001",
5309 => "00000001",
5437 => "00000001",
5565 => "00000001",
5693 => "00000001",
5821 => "00000001",
5949 => "00000001",
6077 => "00000001",
6205 => "00000001",
6333 => "00000001",
6461 => "00000001",
6589 => "00000001",
6717 => "00000001",
6845 => "00000001",
6973 => "00000001",
7101 => "00000001",
7229 => "00000001",
7357 => "00000001",
7485 => "00000001",
7613 => "00000001",
7741 => "00000001",
7869 => "00000001",
7997 => "00000001",
8125 => "00000001",
8253 => "00000001",
8381 => "00000001",
8509 => "00000001",
8637 => "00000001",
8765 => "00000001",
8893 => "00000001",
9021 => "00000001",
9149 => "00000001",
9277 => "00000001",
9405 => "00000001",
9533 => "00000001",
9661 => "00000001",
9789 => "00000001",
9917 => "00000001",
10045 => "00000001",
10173 => "00000001",
10301 => "00000001",
10429 => "00000001",
10557 => "00000001",
10685 => "00000001",
10813 => "00000001",
10941 => "00000001",
11069 => "00000001",
11197 => "00000001",
11325 => "00000001",
11453 => "00000001",
11581 => "00000001",
11709 => "00000001",
11837 => "00000001",
11965 => "00000001",
12093 => "00000001",
12221 => "00000001",
12349 => "00000001",
12477 => "00000001",
12605 => "00000001",
12733 => "00000001",
12861 => "00000001",
12989 => "00000001",
13117 => "00000001",
13245 => "00000001",
13373 => "00000001",
13501 => "00000001",
13629 => "00000001",
13757 => "00000001",
13885 => "00000001",
14013 => "00000001",
14141 => "00000001",
14269 => "00000001",
14397 => "00000001",
14525 => "00000001",
14653 => "00000001",
14781 => "00000001",
14909 => "00000001",
15037 => "00000001",
15165 => "00000001",
15293 => "00000001",
15421 => "00000001",
15549 => "00000001",
15677 => "00000001",
15805 => "00000001",
15933 => "00000001",
16061 => "00000001",
16189 => "00000001",
16317 => "00000001",
67 => "00000001",
195 => "00000001",
323 => "00000001",
451 => "00000001",
579 => "00000001",
707 => "00000001",
835 => "00000001",
963 => "00000001",
1091 => "00000001",
1219 => "00000001",
1347 => "00000001",
1475 => "00000001",
1603 => "00000001",
1731 => "00000001",
1859 => "00000001",
1987 => "00000001",
2115 => "00000001",
2243 => "00000001",
2371 => "00000001",
2499 => "00000001",
2627 => "00000001",
2755 => "00000001",
2883 => "00000001",
3011 => "00000001",
3139 => "00000001",
3267 => "00000001",
3395 => "00000001",
3523 => "00000001",
3651 => "00000001",
3779 => "00000001",
3907 => "00000001",
4035 => "00000001",
4163 => "00000001",
4291 => "00000001",
4419 => "00000001",
4547 => "00000001",
4675 => "00000001",
4803 => "00000001",
4931 => "00000001",
5059 => "00000001",
5187 => "00000001",
5315 => "00000001",
5443 => "00000001",
5571 => "00000001",
5699 => "00000001",
5827 => "00000001",
5955 => "00000001",
6083 => "00000001",
6211 => "00000001",
6339 => "00000001",
6467 => "00000001",
6595 => "00000001",
6723 => "00000001",
6851 => "00000001",
6979 => "00000001",
7107 => "00000001",
7235 => "00000001",
7363 => "00000001",
7491 => "00000001",
7619 => "00000001",
7747 => "00000001",
7875 => "00000001",
8003 => "00000001",
8131 => "00000001",
8259 => "00000001",
8387 => "00000001",
8515 => "00000001",
8643 => "00000001",
8771 => "00000001",
8899 => "00000001",
9027 => "00000001",
9155 => "00000001",
9283 => "00000001",
9411 => "00000001",
9539 => "00000001",
9667 => "00000001",
9795 => "00000001",
9923 => "00000001",
10051 => "00000001",
10179 => "00000001",
10307 => "00000001",
10435 => "00000001",
10563 => "00000001",
10691 => "00000001",
10819 => "00000001",
10947 => "00000001",
11075 => "00000001",
11203 => "00000001",
11331 => "00000001",
11459 => "00000001",
11587 => "00000001",
11715 => "00000001",
11843 => "00000001",
11971 => "00000001",
12099 => "00000001",
12227 => "00000001",
12355 => "00000001",
12483 => "00000001",
12611 => "00000001",
12739 => "00000001",
12867 => "00000001",
12995 => "00000001",
13123 => "00000001",
13251 => "00000001",
13379 => "00000001",
13507 => "00000001",
13635 => "00000001",
13763 => "00000001",
13891 => "00000001",
14019 => "00000001",
14147 => "00000001",
14275 => "00000001",
14403 => "00000001",
14531 => "00000001",
14659 => "00000001",
14787 => "00000001",
14915 => "00000001",
15043 => "00000001",
15171 => "00000001",
15299 => "00000001",
15427 => "00000001",
15555 => "00000001",
15683 => "00000001",
15811 => "00000001",
15939 => "00000001",
16067 => "00000001",
16195 => "00000001",
16323 => "00000001",
73 => "00000001",
201 => "00000001",
329 => "00000001",
457 => "00000001",
585 => "00000001",
713 => "00000001",
841 => "00000001",
969 => "00000001",
1097 => "00000001",
1225 => "00000001",
1353 => "00000001",
1481 => "00000001",
1609 => "00000001",
1737 => "00000001",
1865 => "00000001",
1993 => "00000001",
2121 => "00000001",
2249 => "00000001",
2377 => "00000001",
2505 => "00000001",
2633 => "00000001",
2761 => "00000001",
2889 => "00000001",
3017 => "00000001",
3145 => "00000001",
3273 => "00000001",
3401 => "00000001",
3529 => "00000001",
3657 => "00000001",
3785 => "00000001",
3913 => "00000001",
4041 => "00000001",
4169 => "00000001",
4297 => "00000001",
4425 => "00000001",
4553 => "00000001",
4681 => "00000001",
4809 => "00000001",
4937 => "00000001",
5065 => "00000001",
5193 => "00000001",
5321 => "00000001",
5449 => "00000001",
5577 => "00000001",
5705 => "00000001",
5833 => "00000001",
5961 => "00000001",
6089 => "00000001",
6217 => "00000001",
6345 => "00000001",
6473 => "00000001",
6601 => "00000001",
6729 => "00000001",
6857 => "00000001",
6985 => "00000001",
7113 => "00000001",
7241 => "00000001",
7369 => "00000001",
7497 => "00000001",
7625 => "00000001",
7753 => "00000001",
7881 => "00000001",
8009 => "00000001",
8137 => "00000001",
8265 => "00000001",
8393 => "00000001",
8521 => "00000001",
8649 => "00000001",
8777 => "00000001",
8905 => "00000001",
9033 => "00000001",
9161 => "00000001",
9289 => "00000001",
9417 => "00000001",
9545 => "00000001",
9673 => "00000001",
9801 => "00000001",
9929 => "00000001",
10057 => "00000001",
10185 => "00000001",
10313 => "00000001",
10441 => "00000001",
10569 => "00000001",
10697 => "00000001",
10825 => "00000001",
10953 => "00000001",
11081 => "00000001",
11209 => "00000001",
11337 => "00000001",
11465 => "00000001",
11593 => "00000001",
11721 => "00000001",
11849 => "00000001",
11977 => "00000001",
12105 => "00000001",
12233 => "00000001",
12361 => "00000001",
12489 => "00000001",
12617 => "00000001",
12745 => "00000001",
12873 => "00000001",
13001 => "00000001",
13129 => "00000001",
13257 => "00000001",
13385 => "00000001",
13513 => "00000001",
13641 => "00000001",
13769 => "00000001",
13897 => "00000001",
14025 => "00000001",
14153 => "00000001",
14281 => "00000001",
14409 => "00000001",
14537 => "00000001",
14665 => "00000001",
14793 => "00000001",
14921 => "00000001",
15049 => "00000001",
15177 => "00000001",
15305 => "00000001",
15433 => "00000001",
15561 => "00000001",
15689 => "00000001",
15817 => "00000001",
15945 => "00000001",
16073 => "00000001",
16201 => "00000001",
16329 => "00000001",
79 => "00000010",
207 => "00000010",
335 => "00000010",
463 => "00000010",
591 => "00000010",
719 => "00000010",
847 => "00000010",
975 => "00000010",
1103 => "00000010",
1231 => "00000010",
1359 => "00000010",
1487 => "00000010",
1615 => "00000010",
1743 => "00000010",
1871 => "00000010",
1999 => "00000010",
2127 => "00000010",
2255 => "00000010",
2383 => "00000010",
2511 => "00000010",
2639 => "00000010",
2767 => "00000010",
2895 => "00000010",
3023 => "00000010",
3151 => "00000010",
3279 => "00000010",
3407 => "00000010",
3535 => "00000010",
3663 => "00000010",
3791 => "00000010",
3919 => "00000010",
4047 => "00000010",
4175 => "00000010",
4303 => "00000010",
4431 => "00000010",
4559 => "00000010",
4687 => "00000010",
4815 => "00000010",
4943 => "00000010",
5071 => "00000010",
5199 => "00000010",
5327 => "00000010",
5455 => "00000010",
5583 => "00000010",
5711 => "00000010",
5839 => "00000010",
5967 => "00000010",
6095 => "00000010",
6223 => "00000010",
6351 => "00000010",
6479 => "00000010",
6607 => "00000010",
6735 => "00000010",
6863 => "00000010",
6991 => "00000010",
7119 => "00000010",
7247 => "00000010",
7375 => "00000010",
7503 => "00000010",
7631 => "00000010",
7759 => "00000010",
7887 => "00000010",
8015 => "00000010",
8143 => "00000010",
8271 => "00000010",
8399 => "00000010",
8527 => "00000010",
8655 => "00000010",
8783 => "00000010",
8911 => "00000010",
9039 => "00000010",
9167 => "00000010",
9295 => "00000010",
9423 => "00000010",
9551 => "00000010",
9679 => "00000010",
9807 => "00000010",
9935 => "00000010",
10063 => "00000010",
10191 => "00000010",
10319 => "00000010",
10447 => "00000010",
10575 => "00000010",
10703 => "00000010",
10831 => "00000010",
10959 => "00000010",
11087 => "00000010",
11215 => "00000010",
11343 => "00000010",
11471 => "00000010",
11599 => "00000010",
11727 => "00000010",
11855 => "00000010",
11983 => "00000010",
12111 => "00000010",
12239 => "00000010",
12367 => "00000010",
12495 => "00000010",
12623 => "00000010",
12751 => "00000010",
12879 => "00000010",
13007 => "00000010",
13135 => "00000010",
13263 => "00000010",
13391 => "00000010",
13519 => "00000010",
13647 => "00000010",
13775 => "00000010",
13903 => "00000010",
14031 => "00000010",
14159 => "00000010",
14287 => "00000010",
14415 => "00000010",
14543 => "00000010",
14671 => "00000010",
14799 => "00000010",
14927 => "00000010",
15055 => "00000010",
15183 => "00000010",
15311 => "00000010",
15439 => "00000010",
15567 => "00000010",
15695 => "00000010",
15823 => "00000010",
15951 => "00000010",
16079 => "00000010",
16207 => "00000010",
16335 => "00000010",
    others => (others => '0')
    );

    attribute ram_style : string;
    attribute ram_style of tile_data_map : signal is "block";
    

begin
    -- Write process
    process(i_clk)
        variable write_index : std_logic_vector(13 downto 0);
        variable new_data    : std_logic_vector(7 downto 0);
        variable tile_data : std_logic_vector (7 downto 0);
        variable s_view_index : std_logic_vector (13 downto 0);
    begin
        if rising_edge(i_clk) then
            if (i_ch_we_tileBack = '1') then
                write_index := i_row & i_col;
                --new_data := tile_data_map(to_integer(unsigned(write_index)));
                new_data := (others => '0');
                new_data(4 downto 0) := i_tile_id;
                new_data(5) := i_flip_y;
                new_data(6) := '0';
                new_data(7) := '0';

                -- Update tile_id if required
--                if i_ch_tile_id = '1' then
--                    new_data(4 downto 0) := i_tile_id;
--                end if;

--                -- Update flip_y if required
--                if i_ch_flip_y = '1' then
--                    new_data(5) := i_flip_y;
--                end if;

                -- Write back to BRAM
                tile_data_map(to_integer(unsigned(write_index))) <= new_data;
            end if;
            s_view_index := i_view_y(9 downto 3) & i_view_x(9 downto 3);
            tile_data := tile_data_map(to_integer(unsigned(s_view_index)));
            o_tile_id <= tile_data(4 downto 0);
            o_flip_y  <= tile_data(5);
            o_pix_x   <= i_view_x(2 downto 0);
            o_pix_y   <= i_view_y(2 downto 0);
        end if;
    end process;

end Behavioral;