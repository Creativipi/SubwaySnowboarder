library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity TuileBuffActor is
    Port(
    i_x : in STD_LOGIC_VECTOR (3 downto 0);
    i_y : in STD_LOGIC_VECTOR (3 downto 0);
    i_tile_id : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_x : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_y : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_cc : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_we : in std_logic;
    i_clk : in STD_LOGIC;
    i_tile_id_write : in STD_LOGIC_VECTOR (3 downto 0);
    o_colorCode : out STD_LOGIC_VECTOR (3 downto 0));
end TuileBuffActor;

architecture Behavioral of TuileBuffActor is
constant wh : std_logic_vector (3 downto 0) := "0000"; -- White
constant bl : std_logic_vector (3 downto 0) := "0001"; -- Black
constant ye : std_logic_vector (3 downto 0) := "0010"; -- Yellow
constant dg : std_logic_vector (3 downto 0) := "0011"; -- Dark Green
constant oa : std_logic_vector (3 downto 0) := "0100"; -- Orange
constant bu : std_logic_vector (3 downto 0) := "0101"; -- Blue
constant ge : std_logic_vector (3 downto 0) := "0110"; -- Green
constant lo : std_logic_vector (3 downto 0) := "0111"; -- Light Brown
constant br : std_logic_vector (3 downto 0) := "1000"; -- Brown
constant lg : std_logic_vector (3 downto 0) := "1001"; -- Light Gray
constant gr : std_logic_vector (3 downto 0) := "1010"; -- Gray
constant lb : std_logic_vector (3 downto 0) := "1011"; -- Light Blue
constant sb : std_logic_vector (3 downto 0) := "1100"; -- Sky Blue
constant sa : std_logic_vector (3 downto 0) := "1101"; -- Salmon
constant pi : std_logic_vector (3 downto 0) := "1110"; -- Pink
constant pu : std_logic_vector (3 downto 0) := "1111"; -- Purple

    type tuile_out_array_t is array (0 to 7) of std_logic_vector(3 downto 0);
    signal tuile_outputs : tuile_out_array_t;
    signal tuile_write_enable : std_logic_vector(7 downto 0);
    
    type tile_d_array_t is array (0 to 4095) of std_logic_vector(3 downto 0);
    signal tile_data_map_d : tile_d_array_t :=
    (
0 => pu,
1 => pu,
2 => pu,
3 => pu,
4 => pu,
5 => pu,
6 => pu,
7 => pu,
8 => bu,
9 => pu,
10 => pu,
11 => pu,
12 => pu,
13 => pu,
14 => pu,
15 => pu,
16 => pu,
17 => pu,
18 => pu,
19 => pu,
20 => pu,
21 => pu,
22 => pu,
23 => bu,
24 => wh,
25 => pu,
26 => pu,
27 => pu,
28 => pu,
29 => pu,
30 => pu,
31 => pu,
32 => pu,
33 => pu,
34 => bl,
35 => pu,
36 => pu,
37 => pu,
38 => bu,
39 => wh,
40 => wh,
41 => pu,
42 => pu,
43 => pu,
44 => pu,
45 => pu,
46 => pu,
47 => pu,
48 => pu,
49 => bl,
50 => bl,
51 => bl,
52 => pu,
53 => bu,
54 => wh,
55 => wh,
56 => wh,
57 => pu,
58 => pu,
59 => pu,
60 => pu,
61 => pu,
62 => pu,
63 => pu,
64 => pu,
65 => bl,
66 => bl,
67 => bl,
68 => ye,
69 => wh,
70 => wh,
71 => wh,
72 => wh,
73 => pu,
74 => pu,
75 => pu,
76 => pu,
77 => pu,
78 => pu,
79 => pu,
80 => pu,
81 => pu,
82 => bl,
83 => ye,
84 => bl,
85 => wh,
86 => wh,
87 => wh,
88 => wh,
89 => pu,
90 => pu,
91 => pu,
92 => pu,
93 => pu,
94 => pu,
95 => pu,
96 => pu,
97 => pu,
98 => ye,
99 => bl,
100 => bl,
101 => bl,
102 => wh,
103 => wh,
104 => wh,
105 => pu,
106 => pu,
107 => pu,
108 => pu,
109 => pu,
110 => pu,
111 => pu,
112 => pu,
113 => bu,
114 => wh,
115 => bl,
116 => bl,
117 => bl,
118 => bl,
119 => wh,
120 => bl,
121 => bl,
122 => bl,
123 => bl,
124 => bl,
125 => bl,
126 => pu,
127 => bu,
128 => pu,
129 => bu,
130 => wh,
131 => wh,
132 => bl,
133 => bl,
134 => bl,
135 => bl,
136 => bl,
137 => bl,
138 => bl,
139 => bl,
140 => bl,
141 => bl,
142 => bu,
143 => pu,
144 => bu,
145 => wh,
146 => wh,
147 => wh,
148 => wh,
149 => bl,
150 => bl,
151 => bl,
152 => bl,
153 => bl,
154 => bl,
155 => bl,
156 => bl,
157 => bu,
158 => pu,
159 => pu,
160 => bu,
161 => wh,
162 => wh,
163 => wh,
164 => wh,
165 => wh,
166 => bl,
167 => bl,
168 => bl,
169 => bl,
170 => bl,
171 => bl,
172 => bu,
173 => pu,
174 => pu,
175 => pu,
176 => bu,
177 => wh,
178 => wh,
179 => wh,
180 => wh,
181 => wh,
182 => wh,
183 => bl,
184 => bl,
185 => bl,
186 => wh,
187 => bu,
188 => pu,
189 => pu,
190 => pu,
191 => pu,
192 => bu,
193 => wh,
194 => wh,
195 => wh,
196 => wh,
197 => wh,
198 => wh,
199 => wh,
200 => wh,
201 => wh,
202 => bu,
203 => pu,
204 => pu,
205 => pu,
206 => pu,
207 => pu,
208 => pu,
209 => bu,
210 => wh,
211 => wh,
212 => wh,
213 => wh,
214 => wh,
215 => wh,
216 => wh,
217 => bu,
218 => pu,
219 => pu,
220 => pu,
221 => pu,
222 => pu,
223 => pu,
224 => pu,
225 => pu,
226 => bu,
227 => wh,
228 => wh,
229 => wh,
230 => wh,
231 => bu,
232 => bu,
233 => pu,
234 => pu,
235 => pu,
236 => pu,
237 => pu,
238 => pu,
239 => pu,
240 => pu,
241 => pu,
242 => pu,
243 => bu,
244 => bu,
245 => bu,
246 => bu,
247 => pu,
248 => pu,
249 => pu,
250 => pu,
251 => pu,
252 => pu,
253 => pu,
254 => pu,
255 => pu,
256 => pu,
257 => pu,
258 => pu,
259 => pu,
260 => pu,
261 => pu,
262 => pu,
263 => pu,
264 => pu,
265 => bu,
266 => bu,
267 => bu,
268 => bu,
269 => pu,
270 => pu,
271 => bl,
272 => pu,
273 => pu,
274 => pu,
275 => pu,
276 => pu,
277 => pu,
278 => pu,
279 => bu,
280 => bu,
281 => wh,
282 => wh,
283 => wh,
284 => wh,
285 => bu,
286 => bl,
287 => bl,
288 => pu,
289 => pu,
290 => pu,
291 => pu,
292 => pu,
293 => pu,
294 => bu,
295 => wh,
296 => wh,
297 => wh,
298 => wh,
299 => wh,
300 => wh,
301 => ye,
302 => bl,
303 => bl,
304 => pu,
305 => pu,
306 => pu,
307 => pu,
308 => pu,
309 => bu,
310 => wh,
311 => wh,
312 => wh,
313 => wh,
314 => wh,
315 => wh,
316 => wh,
317 => bl,
318 => ye,
319 => bl,
320 => pu,
321 => pu,
322 => pu,
323 => pu,
324 => bu,
325 => wh,
326 => wh,
327 => wh,
328 => wh,
329 => wh,
330 => wh,
331 => wh,
332 => bl,
333 => bl,
334 => bl,
335 => bu,
336 => pu,
337 => pu,
338 => pu,
339 => bu,
340 => wh,
341 => wh,
342 => wh,
343 => wh,
344 => wh,
345 => wh,
346 => wh,
347 => bl,
348 => bl,
349 => bl,
350 => wh,
351 => bu,
352 => pu,
353 => pu,
354 => bu,
355 => wh,
356 => wh,
357 => wh,
358 => wh,
359 => wh,
360 => wh,
361 => bl,
362 => bl,
363 => bl,
364 => bl,
365 => bl,
366 => wh,
367 => bu,
368 => pu,
369 => bu,
370 => wh,
371 => wh,
372 => wh,
373 => wh,
374 => wh,
375 => bl,
376 => bl,
377 => bl,
378 => bl,
379 => bl,
380 => bl,
381 => wh,
382 => wh,
383 => bu,
384 => bu,
385 => wh,
386 => ye,
387 => ye,
388 => ye,
389 => ye,
390 => bl,
391 => bl,
392 => bl,
393 => bl,
394 => bl,
395 => bl,
396 => wh,
397 => wh,
398 => bu,
399 => pu,
400 => wh,
401 => ye,
402 => bl,
403 => bl,
404 => bl,
405 => bl,
406 => ye,
407 => bl,
408 => bl,
409 => bl,
410 => bl,
411 => wh,
412 => wh,
413 => bu,
414 => pu,
415 => pu,
416 => ye,
417 => bl,
418 => bl,
419 => bl,
420 => bl,
421 => bl,
422 => bl,
423 => ye,
424 => bl,
425 => bl,
426 => bl,
427 => wh,
428 => bu,
429 => pu,
430 => pu,
431 => pu,
432 => ye,
433 => bl,
434 => bl,
435 => bl,
436 => bl,
437 => bl,
438 => bl,
439 => ye,
440 => bl,
441 => bl,
442 => wh,
443 => bu,
444 => pu,
445 => pu,
446 => pu,
447 => pu,
448 => ye,
449 => bl,
450 => bl,
451 => bl,
452 => bl,
453 => bl,
454 => bl,
455 => ye,
456 => bl,
457 => wh,
458 => bu,
459 => pu,
460 => pu,
461 => pu,
462 => pu,
463 => pu,
464 => ye,
465 => bl,
466 => bl,
467 => bl,
468 => bl,
469 => bl,
470 => bl,
471 => ye,
472 => wh,
473 => bu,
474 => pu,
475 => pu,
476 => pu,
477 => pu,
478 => pu,
479 => pu,
480 => bl,
481 => ye,
482 => bl,
483 => bl,
484 => bl,
485 => bl,
486 => ye,
487 => wh,
488 => bu,
489 => pu,
490 => pu,
491 => pu,
492 => pu,
493 => pu,
494 => pu,
495 => pu,
496 => bl,
497 => bl,
498 => ye,
499 => ye,
500 => ye,
501 => ye,
502 => wh,
503 => bu,
504 => pu,
505 => pu,
506 => pu,
507 => pu,
508 => pu,
509 => pu,
510 => pu,
511 => pu,
512 => pu,
513 => pu,
514 => pu,
515 => pu,
516 => pu,
517 => pu,
518 => pu,
519 => bl,
520 => bl,
521 => pu,
522 => pu,
523 => pu,
524 => pu,
525 => pu,
526 => pu,
527 => pu,
528 => pu,
529 => pu,
530 => pu,
531 => pu,
532 => pu,
533 => pu,
534 => pu,
535 => bl,
536 => bl,
537 => bl,
538 => pu,
539 => pu,
540 => pu,
541 => pu,
542 => pu,
543 => pu,
544 => pu,
545 => pu,
546 => pu,
547 => pu,
548 => pu,
549 => pu,
550 => bu,
551 => bl,
552 => bl,
553 => bl,
554 => bu,
555 => pu,
556 => pu,
557 => pu,
558 => pu,
559 => pu,
560 => pu,
561 => pu,
562 => pu,
563 => pu,
564 => pu,
565 => bu,
566 => wh,
567 => wh,
568 => ye,
569 => ye,
570 => wh,
571 => bu,
572 => pu,
573 => pu,
574 => pu,
575 => pu,
576 => pu,
577 => pu,
578 => pu,
579 => pu,
580 => bu,
581 => wh,
582 => wh,
583 => wh,
584 => bl,
585 => bl,
586 => wh,
587 => wh,
588 => bu,
589 => pu,
590 => pu,
591 => pu,
592 => pu,
593 => pu,
594 => pu,
595 => pu,
596 => bu,
597 => wh,
598 => wh,
599 => wh,
600 => bl,
601 => bl,
602 => bl,
603 => wh,
604 => bu,
605 => pu,
606 => pu,
607 => pu,
608 => pu,
609 => pu,
610 => pu,
611 => bu,
612 => wh,
613 => wh,
614 => wh,
615 => wh,
616 => bl,
617 => bl,
618 => bl,
619 => wh,
620 => wh,
621 => bu,
622 => pu,
623 => pu,
624 => pu,
625 => pu,
626 => pu,
627 => bu,
628 => wh,
629 => wh,
630 => wh,
631 => wh,
632 => bl,
633 => bl,
634 => bl,
635 => wh,
636 => wh,
637 => bu,
638 => pu,
639 => pu,
640 => pu,
641 => pu,
642 => pu,
643 => bu,
644 => wh,
645 => wh,
646 => wh,
647 => bl,
648 => bl,
649 => bl,
650 => bl,
651 => wh,
652 => wh,
653 => bu,
654 => pu,
655 => pu,
656 => pu,
657 => pu,
658 => pu,
659 => bu,
660 => wh,
661 => wh,
662 => wh,
663 => bl,
664 => bl,
665 => bl,
666 => bl,
667 => wh,
668 => wh,
669 => bu,
670 => pu,
671 => pu,
672 => pu,
673 => pu,
674 => pu,
675 => bu,
676 => wh,
677 => wh,
678 => bl,
679 => bl,
680 => bl,
681 => bl,
682 => bl,
683 => bl,
684 => wh,
685 => bu,
686 => pu,
687 => pu,
688 => pu,
689 => pu,
690 => pu,
691 => bu,
692 => wh,
693 => wh,
694 => bl,
695 => bl,
696 => bl,
697 => bl,
698 => bl,
699 => bl,
700 => wh,
701 => bu,
702 => pu,
703 => pu,
704 => pu,
705 => pu,
706 => pu,
707 => bu,
708 => wh,
709 => wh,
710 => ye,
711 => ye,
712 => ye,
713 => ye,
714 => bl,
715 => bl,
716 => wh,
717 => bu,
718 => pu,
719 => pu,
720 => pu,
721 => pu,
722 => pu,
723 => bu,
724 => wh,
725 => ye,
726 => bl,
727 => bl,
728 => bl,
729 => bl,
730 => ye,
731 => bl,
732 => wh,
733 => bu,
734 => pu,
735 => pu,
736 => pu,
737 => pu,
738 => pu,
739 => bu,
740 => ye,
741 => bl,
742 => bl,
743 => bl,
744 => bl,
745 => bl,
746 => bl,
747 => ye,
748 => wh,
749 => bu,
750 => pu,
751 => pu,
752 => pu,
753 => pu,
754 => pu,
755 => bu,
756 => ye,
757 => bl,
758 => bl,
759 => bl,
760 => bl,
761 => bl,
762 => bl,
763 => ye,
764 => wh,
765 => bu,
766 => pu,
767 => pu,
768 => pu,
769 => pu,
770 => pu,
771 => bu,
772 => ye,
773 => bl,
774 => bl,
775 => bl,
776 => bl,
777 => bl,
778 => bl,
779 => ye,
780 => wh,
781 => bu,
782 => pu,
783 => pu,
784 => pu,
785 => pu,
786 => pu,
787 => bu,
788 => ye,
789 => bl,
790 => bl,
791 => bl,
792 => bl,
793 => bl,
794 => bl,
795 => ye,
796 => wh,
797 => bu,
798 => pu,
799 => pu,
800 => pu,
801 => pu,
802 => pu,
803 => bu,
804 => wh,
805 => ye,
806 => bl,
807 => bl,
808 => bl,
809 => bl,
810 => ye,
811 => bl,
812 => wh,
813 => bu,
814 => pu,
815 => pu,
816 => pu,
817 => pu,
818 => pu,
819 => bu,
820 => wh,
821 => wh,
822 => ye,
823 => ye,
824 => ye,
825 => ye,
826 => bl,
827 => bl,
828 => wh,
829 => bu,
830 => pu,
831 => pu,
832 => pu,
833 => pu,
834 => pu,
835 => bu,
836 => wh,
837 => wh,
838 => wh,
839 => bl,
840 => bl,
841 => bl,
842 => bl,
843 => bl,
844 => wh,
845 => bu,
846 => pu,
847 => pu,
848 => pu,
849 => pu,
850 => pu,
851 => bu,
852 => wh,
853 => wh,
854 => wh,
855 => bl,
856 => bl,
857 => bl,
858 => bl,
859 => bl,
860 => wh,
861 => bu,
862 => pu,
863 => pu,
864 => pu,
865 => pu,
866 => pu,
867 => bu,
868 => wh,
869 => wh,
870 => wh,
871 => bl,
872 => bl,
873 => bl,
874 => bl,
875 => wh,
876 => wh,
877 => bu,
878 => pu,
879 => pu,
880 => pu,
881 => pu,
882 => pu,
883 => bu,
884 => wh,
885 => wh,
886 => wh,
887 => bl,
888 => bl,
889 => bl,
890 => bl,
891 => wh,
892 => wh,
893 => bu,
894 => pu,
895 => pu,
896 => pu,
897 => pu,
898 => pu,
899 => bu,
900 => wh,
901 => wh,
902 => bl,
903 => bl,
904 => bl,
905 => bl,
906 => wh,
907 => wh,
908 => wh,
909 => bu,
910 => pu,
911 => pu,
912 => pu,
913 => pu,
914 => pu,
915 => bu,
916 => wh,
917 => wh,
918 => bl,
919 => bl,
920 => bl,
921 => bl,
922 => wh,
923 => wh,
924 => wh,
925 => bu,
926 => pu,
927 => pu,
928 => pu,
929 => pu,
930 => pu,
931 => bu,
932 => wh,
933 => bl,
934 => bl,
935 => bl,
936 => bl,
937 => wh,
938 => wh,
939 => wh,
940 => wh,
941 => bu,
942 => pu,
943 => pu,
944 => pu,
945 => pu,
946 => pu,
947 => bu,
948 => bl,
949 => ye,
950 => bl,
951 => bl,
952 => wh,
953 => wh,
954 => wh,
955 => wh,
956 => wh,
957 => bu,
958 => pu,
959 => pu,
960 => pu,
961 => pu,
962 => bl,
963 => bl,
964 => bl,
965 => ye,
966 => bl,
967 => wh,
968 => wh,
969 => wh,
970 => wh,
971 => wh,
972 => bu,
973 => pu,
974 => pu,
975 => pu,
976 => pu,
977 => pu,
978 => bl,
979 => bl,
980 => bl,
981 => wh,
982 => wh,
983 => wh,
984 => wh,
985 => wh,
986 => wh,
987 => wh,
988 => bu,
989 => pu,
990 => pu,
991 => pu,
992 => pu,
993 => pu,
994 => pu,
995 => pu,
996 => pu,
997 => bu,
998 => wh,
999 => wh,
1000 => wh,
1001 => wh,
1002 => wh,
1003 => bu,
1004 => pu,
1005 => pu,
1006 => pu,
1007 => pu,
1008 => pu,
1009 => pu,
1010 => pu,
1011 => pu,
1012 => pu,
1013 => pu,
1014 => bu,
1015 => bu,
1016 => bu,
1017 => bu,
1018 => bu,
1019 => pu,
1020 => pu,
1021 => pu,
1022 => pu,
1023 => pu,
1024 => pu,
1025 => pu,
1026 => pu,
1027 => pu,
1028 => pu,
1029 => pu,
1030 => pu,
1031 => pu,
1032 => pu,
1033 => pu,
1034 => pu,
1035 => pu,
1036 => pu,
1037 => pu,
1038 => pu,
1039 => pu,
1040 => pu,
1041 => pu,
1042 => pu,
1043 => bl,
1044 => bl,
1045 => bl,
1046 => pu,
1047 => pu,
1048 => pu,
1049 => pu,
1050 => pu,
1051 => pu,
1052 => pu,
1053 => pu,
1054 => pu,
1055 => pu,
1056 => pu,
1057 => pu,
1058 => bl,
1059 => wh,
1060 => ye,
1061 => ye,
1062 => bl,
1063 => pu,
1064 => pu,
1065 => pu,
1066 => pu,
1067 => pu,
1068 => pu,
1069 => pu,
1070 => pu,
1071 => pu,
1072 => pu,
1073 => bl,
1074 => lg,
1075 => wh,
1076 => wh,
1077 => lg,
1078 => gr,
1079 => bl,
1080 => bl,
1081 => pu,
1082 => pu,
1083 => pu,
1084 => pu,
1085 => pu,
1086 => pu,
1087 => pu,
1088 => bl,
1089 => wh,
1090 => wh,
1091 => wh,
1092 => wh,
1093 => wh,
1094 => wh,
1095 => wh,
1096 => lg,
1097 => bl,
1098 => pu,
1099 => pu,
1100 => pu,
1101 => pu,
1102 => pu,
1103 => pu,
1104 => bl,
1105 => ge,
1106 => wh,
1107 => ye,
1108 => ye,
1109 => ye,
1110 => ye,
1111 => ye,
1112 => wh,
1113 => ge,
1114 => bl,
1115 => bl,
1116 => pu,
1117 => pu,
1118 => pu,
1119 => pu,
1120 => bl,
1121 => ge,
1122 => wh,
1123 => lg,
1124 => ye,
1125 => oa,
1126 => ye,
1127 => oa,
1128 => wh,
1129 => ge,
1130 => ge,
1131 => ge,
1132 => bl,
1133 => pu,
1134 => pu,
1135 => pu,
1136 => pu,
1137 => bl,
1138 => lg,
1139 => oa,
1140 => ye,
1141 => ye,
1142 => oa,
1143 => ye,
1144 => lg,
1145 => dg,
1146 => dg,
1147 => ge,
1148 => dg,
1149 => bl,
1150 => pu,
1151 => pu,
1152 => pu,
1153 => pu,
1154 => bl,
1155 => oa,
1156 => oa,
1157 => oa,
1158 => lg,
1159 => oa,
1160 => wh,
1161 => wh,
1162 => wh,
1163 => wh,
1164 => wh,
1165 => wh,
1166 => bl,
1167 => pu,
1168 => pu,
1169 => pu,
1170 => pu,
1171 => bl,
1172 => oa,
1173 => oa,
1174 => wh,
1175 => wh,
1176 => wh,
1177 => ge,
1178 => ge,
1179 => ge,
1180 => wh,
1181 => oa,
1182 => oa,
1183 => bl,
1184 => pu,
1185 => pu,
1186 => pu,
1187 => pu,
1188 => bl,
1189 => wh,
1190 => wh,
1191 => wh,
1192 => dg,
1193 => ge,
1194 => dg,
1195 => dg,
1196 => dg,
1197 => wh,
1198 => oa,
1199 => bl,
1200 => pu,
1201 => pu,
1202 => pu,
1203 => pu,
1204 => pu,
1205 => bl,
1206 => wh,
1207 => wh,
1208 => wh,
1209 => wh,
1210 => wh,
1211 => dg,
1212 => dg,
1213 => wh,
1214 => wh,
1215 => bl,
1216 => pu,
1217 => pu,
1218 => pu,
1219 => pu,
1220 => pu,
1221 => pu,
1222 => bl,
1223 => lg,
1224 => gr,
1225 => wh,
1226 => wh,
1227 => dg,
1228 => dg,
1229 => wh,
1230 => bl,
1231 => pu,
1232 => pu,
1233 => pu,
1234 => pu,
1235 => pu,
1236 => pu,
1237 => pu,
1238 => pu,
1239 => bl,
1240 => bl,
1241 => gr,
1242 => ge,
1243 => dg,
1244 => wh,
1245 => lg,
1246 => bl,
1247 => pu,
1248 => pu,
1249 => pu,
1250 => pu,
1251 => pu,
1252 => pu,
1253 => pu,
1254 => pu,
1255 => pu,
1256 => pu,
1257 => bl,
1258 => bl,
1259 => lg,
1260 => wh,
1261 => bl,
1262 => pu,
1263 => pu,
1264 => pu,
1265 => pu,
1266 => pu,
1267 => pu,
1268 => pu,
1269 => pu,
1270 => pu,
1271 => pu,
1272 => pu,
1273 => pu,
1274 => pu,
1275 => bl,
1276 => bl,
1277 => pu,
1278 => pu,
1279 => pu,
1280 => pu,
1281 => pu,
1282 => pu,
1283 => pu,
1284 => pu,
1285 => pu,
1286 => pu,
1287 => pu,
1288 => pu,
1289 => pu,
1290 => pu,
1291 => pu,
1292 => pu,
1293 => pu,
1294 => pu,
1295 => pu,
1296 => pu,
1297 => pu,
1298 => pu,
1299 => pu,
1300 => pu,
1301 => bl,
1302 => bl,
1303 => bl,
1304 => bl,
1305 => bl,
1306 => bl,
1307 => pu,
1308 => pu,
1309 => pu,
1310 => pu,
1311 => pu,
1312 => pu,
1313 => pu,
1314 => pu,
1315 => pu,
1316 => bl,
1317 => ge,
1318 => wh,
1319 => lg,
1320 => wh,
1321 => wh,
1322 => ye,
1323 => bl,
1324 => pu,
1325 => pu,
1326 => pu,
1327 => pu,
1328 => pu,
1329 => pu,
1330 => pu,
1331 => bl,
1332 => ge,
1333 => wh,
1334 => wh,
1335 => ye,
1336 => wh,
1337 => wh,
1338 => lg,
1339 => ye,
1340 => bl,
1341 => pu,
1342 => pu,
1343 => pu,
1344 => pu,
1345 => pu,
1346 => pu,
1347 => bl,
1348 => wh,
1349 => wh,
1350 => wh,
1351 => ye,
1352 => ye,
1353 => wh,
1354 => wh,
1355 => gr,
1356 => bl,
1357 => pu,
1358 => pu,
1359 => pu,
1360 => pu,
1361 => pu,
1362 => pu,
1363 => bl,
1364 => oa,
1365 => oa,
1366 => ye,
1367 => oa,
1368 => ye,
1369 => ye,
1370 => wh,
1371 => lg,
1372 => bl,
1373 => pu,
1374 => pu,
1375 => pu,
1376 => pu,
1377 => pu,
1378 => pu,
1379 => bl,
1380 => oa,
1381 => oa,
1382 => oa,
1383 => ye,
1384 => ye,
1385 => ye,
1386 => wh,
1387 => ge,
1388 => bl,
1389 => pu,
1390 => pu,
1391 => pu,
1392 => pu,
1393 => pu,
1394 => pu,
1395 => bl,
1396 => oa,
1397 => oa,
1398 => ye,
1399 => oa,
1400 => ye,
1401 => wh,
1402 => ge,
1403 => ge,
1404 => bl,
1405 => pu,
1406 => pu,
1407 => pu,
1408 => pu,
1409 => pu,
1410 => pu,
1411 => bl,
1412 => wh,
1413 => wh,
1414 => wh,
1415 => wh,
1416 => wh,
1417 => ge,
1418 => ge,
1419 => ge,
1420 => bl,
1421 => pu,
1422 => pu,
1423 => pu,
1424 => pu,
1425 => pu,
1426 => pu,
1427 => bl,
1428 => wh,
1429 => wh,
1430 => ge,
1431 => ge,
1432 => wh,
1433 => wh,
1434 => dg,
1435 => dg,
1436 => bl,
1437 => pu,
1438 => pu,
1439 => pu,
1440 => pu,
1441 => pu,
1442 => pu,
1443 => bl,
1444 => lg,
1445 => ge,
1446 => wh,
1447 => ge,
1448 => ge,
1449 => wh,
1450 => wh,
1451 => dg,
1452 => bl,
1453 => pu,
1454 => pu,
1455 => pu,
1456 => pu,
1457 => pu,
1458 => pu,
1459 => bl,
1460 => gr,
1461 => wh,
1462 => wh,
1463 => dg,
1464 => ge,
1465 => wh,
1466 => wh,
1467 => wh,
1468 => bl,
1469 => pu,
1470 => pu,
1471 => pu,
1472 => pu,
1473 => pu,
1474 => pu,
1475 => bl,
1476 => lg,
1477 => dg,
1478 => dg,
1479 => dg,
1480 => dg,
1481 => wh,
1482 => oa,
1483 => oa,
1484 => bl,
1485 => pu,
1486 => pu,
1487 => pu,
1488 => pu,
1489 => pu,
1490 => pu,
1491 => pu,
1492 => bl,
1493 => lg,
1494 => dg,
1495 => dg,
1496 => lg,
1497 => wh,
1498 => oa,
1499 => bl,
1500 => pu,
1501 => pu,
1502 => pu,
1503 => pu,
1504 => pu,
1505 => pu,
1506 => pu,
1507 => pu,
1508 => pu,
1509 => bl,
1510 => bl,
1511 => bl,
1512 => bl,
1513 => bl,
1514 => bl,
1515 => pu,
1516 => pu,
1517 => pu,
1518 => pu,
1519 => pu,
1520 => pu,
1521 => pu,
1522 => pu,
1523 => pu,
1524 => pu,
1525 => pu,
1526 => pu,
1527 => pu,
1528 => pu,
1529 => pu,
1530 => pu,
1531 => pu,
1532 => pu,
1533 => pu,
1534 => pu,
1535 => pu,
1536 => pu,
1537 => pu,
1538 => pu,
1539 => pu,
1540 => pu,
1541 => pu,
1542 => pu,
1543 => pu,
1544 => pu,
1545 => pu,
1546 => pu,
1547 => pu,
1548 => pu,
1549 => pu,
1550 => pu,
1551 => pu,
1552 => pu,
1553 => pu,
1554 => pu,
1555 => pu,
1556 => pu,
1557 => pu,
1558 => pu,
1559 => pu,
1560 => pu,
1561 => pu,
1562 => pu,
1563 => bl,
1564 => bl,
1565 => pu,
1566 => pu,
1567 => pu,
1568 => pu,
1569 => pu,
1570 => pu,
1571 => pu,
1572 => pu,
1573 => pu,
1574 => pu,
1575 => pu,
1576 => pu,
1577 => pu,
1578 => bl,
1579 => ge,
1580 => ge,
1581 => bl,
1582 => pu,
1583 => pu,
1584 => pu,
1585 => pu,
1586 => pu,
1587 => pu,
1588 => pu,
1589 => pu,
1590 => pu,
1591 => pu,
1592 => bl,
1593 => bl,
1594 => wh,
1595 => wh,
1596 => wh,
1597 => wh,
1598 => bl,
1599 => pu,
1600 => pu,
1601 => pu,
1602 => pu,
1603 => pu,
1604 => pu,
1605 => pu,
1606 => bl,
1607 => bl,
1608 => oa,
1609 => oa,
1610 => oa,
1611 => ye,
1612 => ye,
1613 => wh,
1614 => lg,
1615 => bl,
1616 => pu,
1617 => pu,
1618 => pu,
1619 => pu,
1620 => pu,
1621 => bl,
1622 => wh,
1623 => oa,
1624 => oa,
1625 => ye,
1626 => ye,
1627 => ye,
1628 => ye,
1629 => wh,
1630 => wh,
1631 => bl,
1632 => pu,
1633 => pu,
1634 => pu,
1635 => bl,
1636 => bl,
1637 => wh,
1638 => wh,
1639 => wh,
1640 => oa,
1641 => oa,
1642 => oa,
1643 => ye,
1644 => ye,
1645 => wh,
1646 => ye,
1647 => bl,
1648 => pu,
1649 => pu,
1650 => bl,
1651 => wh,
1652 => lg,
1653 => ge,
1654 => wh,
1655 => wh,
1656 => lg,
1657 => oa,
1658 => ye,
1659 => ye,
1660 => wh,
1661 => lg,
1662 => ye,
1663 => bl,
1664 => pu,
1665 => bl,
1666 => gr,
1667 => lg,
1668 => wh,
1669 => dg,
1670 => ge,
1671 => wh,
1672 => oa,
1673 => ye,
1674 => oa,
1675 => ye,
1676 => wh,
1677 => gr,
1678 => bl,
1679 => pu,
1680 => bl,
1681 => lg,
1682 => dg,
1683 => wh,
1684 => wh,
1685 => ge,
1686 => dg,
1687 => wh,
1688 => wh,
1689 => wh,
1690 => wh,
1691 => wh,
1692 => wh,
1693 => bl,
1694 => pu,
1695 => pu,
1696 => bl,
1697 => lg,
1698 => dg,
1699 => ge,
1700 => ge,
1701 => dg,
1702 => ge,
1703 => wh,
1704 => dg,
1705 => ge,
1706 => ge,
1707 => lg,
1708 => bl,
1709 => pu,
1710 => pu,
1711 => pu,
1712 => bl,
1713 => wh,
1714 => wh,
1715 => dg,
1716 => dg,
1717 => ge,
1718 => wh,
1719 => wh,
1720 => ge,
1721 => dg,
1722 => bl,
1723 => bl,
1724 => pu,
1725 => pu,
1726 => pu,
1727 => pu,
1728 => pu,
1729 => bl,
1730 => lg,
1731 => wh,
1732 => wh,
1733 => wh,
1734 => wh,
1735 => wh,
1736 => dg,
1737 => bl,
1738 => pu,
1739 => pu,
1740 => pu,
1741 => pu,
1742 => pu,
1743 => pu,
1744 => pu,
1745 => pu,
1746 => bl,
1747 => wh,
1748 => wh,
1749 => oa,
1750 => wh,
1751 => dg,
1752 => bl,
1753 => pu,
1754 => pu,
1755 => pu,
1756 => pu,
1757 => pu,
1758 => pu,
1759 => pu,
1760 => pu,
1761 => pu,
1762 => pu,
1763 => bl,
1764 => oa,
1765 => oa,
1766 => bl,
1767 => bl,
1768 => pu,
1769 => pu,
1770 => pu,
1771 => pu,
1772 => pu,
1773 => pu,
1774 => pu,
1775 => pu,
1776 => pu,
1777 => pu,
1778 => pu,
1779 => pu,
1780 => bl,
1781 => bl,
1782 => pu,
1783 => pu,
1784 => pu,
1785 => pu,
1786 => pu,
1787 => pu,
1788 => pu,
1789 => pu,
1790 => pu,
1791 => pu,
1792 => pu,
1793 => pu,
1794 => pu,
1795 => pu,
1796 => pu,
1797 => pu,
1798 => pu,
1799 => pu,
1800 => pu,
1801 => pu,
1802 => pu,
1803 => pu,
1804 => pu,
1805 => pu,
1806 => pu,
1807 => pu,
1808 => pu,
1809 => pu,
1810 => pu,
1811 => pu,
1812 => pu,
1813 => pu,
1814 => pu,
1815 => pu,
1816 => pu,
1817 => pu,
1818 => pu,
1819 => pu,
1820 => pu,
1821 => pu,
1822 => pu,
1823 => pu,
1824 => pu,
1825 => pu,
1826 => pu,
1827 => pu,
1828 => pu,
1829 => pu,
1830 => pu,
1831 => pu,
1832 => pu,
1833 => pu,
1834 => pu,
1835 => pu,
1836 => pu,
1837 => pu,
1838 => pu,
1839 => pu,
1840 => pu,
1841 => pu,
1842 => bl,
1843 => bl,
1844 => bl,
1845 => bl,
1846 => bl,
1847 => bl,
1848 => bl,
1849 => bl,
1850 => bl,
1851 => bl,
1852 => bl,
1853 => bl,
1854 => pu,
1855 => pu,
1856 => pu,
1857 => bl,
1858 => ye,
1859 => lg,
1860 => gr,
1861 => wh,
1862 => ge,
1863 => ge,
1864 => dg,
1865 => ge,
1866 => dg,
1867 => wh,
1868 => wh,
1869 => oa,
1870 => bl,
1871 => pu,
1872 => bl,
1873 => ye,
1874 => wh,
1875 => lg,
1876 => wh,
1877 => ye,
1878 => wh,
1879 => ge,
1880 => dg,
1881 => dg,
1882 => wh,
1883 => wh,
1884 => wh,
1885 => oa,
1886 => oa,
1887 => bl,
1888 => bl,
1889 => wh,
1890 => wh,
1891 => wh,
1892 => ye,
1893 => ye,
1894 => ye,
1895 => wh,
1896 => ge,
1897 => wh,
1898 => wh,
1899 => wh,
1900 => wh,
1901 => wh,
1902 => wh,
1903 => bl,
1904 => bl,
1905 => lg,
1906 => wh,
1907 => ye,
1908 => ye,
1909 => oa,
1910 => oa,
1911 => ye,
1912 => wh,
1913 => wh,
1914 => ge,
1915 => ge,
1916 => dg,
1917 => dg,
1918 => wh,
1919 => bl,
1920 => bl,
1921 => wh,
1922 => ye,
1923 => ye,
1924 => oa,
1925 => ye,
1926 => oa,
1927 => ye,
1928 => wh,
1929 => ge,
1930 => dg,
1931 => dg,
1932 => ge,
1933 => dg,
1934 => lg,
1935 => bl,
1936 => bl,
1937 => ge,
1938 => wh,
1939 => wh,
1940 => ye,
1941 => oa,
1942 => oa,
1943 => wh,
1944 => wh,
1945 => ge,
1946 => dg,
1947 => wh,
1948 => wh,
1949 => dg,
1950 => dg,
1951 => bl,
1952 => bl,
1953 => ge,
1954 => wh,
1955 => wh,
1956 => oa,
1957 => oa,
1958 => oa,
1959 => wh,
1960 => wh,
1961 => ge,
1962 => dg,
1963 => wh,
1964 => wh,
1965 => dg,
1966 => dg,
1967 => bl,
1968 => pu,
1969 => bl,
1970 => dg,
1971 => wh,
1972 => oa,
1973 => oa,
1974 => oa,
1975 => wh,
1976 => wh,
1977 => wh,
1978 => dg,
1979 => lg,
1980 => gr,
1981 => lg,
1982 => bl,
1983 => pu,
1984 => pu,
1985 => pu,
1986 => bl,
1987 => bl,
1988 => bl,
1989 => bl,
1990 => bl,
1991 => bl,
1992 => bl,
1993 => bl,
1994 => bl,
1995 => bl,
1996 => bl,
1997 => bl,
1998 => pu,
1999 => pu,
2000 => pu,
2001 => pu,
2002 => pu,
2003 => pu,
2004 => pu,
2005 => pu,
2006 => pu,
2007 => pu,
2008 => pu,
2009 => pu,
2010 => pu,
2011 => pu,
2012 => pu,
2013 => pu,
2014 => pu,
2015 => pu,
2016 => pu,
2017 => pu,
2018 => pu,
2019 => pu,
2020 => pu,
2021 => pu,
2022 => pu,
2023 => pu,
2024 => pu,
2025 => pu,
2026 => pu,
2027 => pu,
2028 => pu,
2029 => pu,
2030 => pu,
2031 => pu,
2032 => pu,
2033 => pu,
2034 => pu,
2035 => pu,
2036 => pu,
2037 => pu,
2038 => pu,
2039 => pu,
2040 => pu,
2041 => pu,
2042 => pu,
2043 => pu,
2044 => pu,
2045 => pu,
2046 => pu,
2047 => pu,
others => pu
    ); 
    
    attribute ram_style : string;
    attribute ram_style of tile_data_map_d : signal is "block";
begin
    
      process(i_tile_id, i_x, i_y)
          variable readIndex : std_logic_vector (11 downto 0);
          variable readIndex_int : integer;
          begin
          readIndex := i_tile_id & i_y & i_x;
          readIndex_int := to_integer(unsigned(readIndex));
          o_colorCode <= tile_data_map_d(readIndex_int);
      end process;
      
      process(i_clk)
      variable writeIndex : std_logic_vector (11 downto 0);
      variable writeIndex_int : integer;
      begin
        if rising_edge(i_clk) then
            if i_ch_we = '1' then
                writeIndex := i_tile_id_write & i_ch_y & i_ch_x;
                writeIndex_int := to_integer(unsigned(writeIndex));
                tile_data_map_d(writeIndex_int) <= i_ch_cc;
            end if;
        end if;
      end process;

end Behavioral;
