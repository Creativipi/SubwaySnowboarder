library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity TuileBuffActor is
    Port(
    i_x : in STD_LOGIC_VECTOR (3 downto 0);
    i_y : in STD_LOGIC_VECTOR (3 downto 0);
    i_tile_id : in STD_LOGIC_VECTOR (2 downto 0);
    i_ch_x : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_y : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_cc : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_we : in std_logic;
    i_clk : in STD_LOGIC;
    i_flip_y : in STD_LOGIC;
    i_tile_id_write : in STD_LOGIC_VECTOR (2 downto 0);
    o_colorCode : out STD_LOGIC_VECTOR (3 downto 0));
end TuileBuffActor;

architecture Behavioral of TuileBuffActor is
constant wh : std_logic_vector (3 downto 0) := "0000"; -- White
constant bl : std_logic_vector (3 downto 0) := "0001"; -- Black
constant ye : std_logic_vector (3 downto 0) := "0010"; -- Yellow
constant dg : std_logic_vector (3 downto 0) := "0011"; -- Dark Green
constant oa : std_logic_vector (3 downto 0) := "0100"; -- Orange
constant bu : std_logic_vector (3 downto 0) := "0101"; -- Blue
constant ge : std_logic_vector (3 downto 0) := "0110"; -- Green
constant lo : std_logic_vector (3 downto 0) := "0111"; -- Light Brown
constant br : std_logic_vector (3 downto 0) := "1000"; -- Brown
constant lg : std_logic_vector (3 downto 0) := "1001"; -- Light Gray
constant gr : std_logic_vector (3 downto 0) := "1010"; -- Gray
constant lb : std_logic_vector (3 downto 0) := "1011"; -- Light Blue
constant sb : std_logic_vector (3 downto 0) := "1100"; -- Sky Blue
constant sa : std_logic_vector (3 downto 0) := "1101"; -- Salmon
constant pi : std_logic_vector (3 downto 0) := "1110"; -- Pink
constant pu : std_logic_vector (3 downto 0) := "1111"; -- Purple

    type tuile_out_array_t is array (0 to 7) of std_logic_vector(3 downto 0);
    signal tuile_outputs : tuile_out_array_t;
    signal tuile_write_enable : std_logic_vector(7 downto 0);
    
    type tile_d_array_t is array (0 to 2047) of std_logic_vector(3 downto 0);
    signal tile_data_map_d : tile_d_array_t :=
    (
0 => wh,
1 => wh,
2 => wh,
3 => wh,
4 => wh,
5 => wh,
6 => wh,
7 => wh,
8 => bu,
9 => wh,
10 => wh,
11 => wh,
12 => wh,
13 => wh,
14 => wh,
15 => wh,
16 => wh,
17 => wh,
18 => wh,
19 => wh,
20 => wh,
21 => wh,
22 => wh,
23 => bu,
24 => wh,
25 => wh,
26 => wh,
27 => wh,
28 => wh,
29 => wh,
30 => wh,
31 => wh,
32 => wh,
33 => wh,
34 => bl,
35 => wh,
36 => wh,
37 => wh,
38 => bu,
39 => wh,
40 => wh,
41 => wh,
42 => wh,
43 => wh,
44 => wh,
45 => wh,
46 => wh,
47 => wh,
48 => wh,
49 => bl,
50 => bl,
51 => bl,
52 => wh,
53 => bu,
54 => wh,
55 => wh,
56 => wh,
57 => wh,
58 => wh,
59 => wh,
60 => wh,
61 => wh,
62 => wh,
63 => wh,
64 => wh,
65 => bl,
66 => bl,
67 => bl,
68 => oa,
69 => wh,
70 => wh,
71 => wh,
72 => wh,
73 => wh,
74 => wh,
75 => wh,
76 => wh,
77 => wh,
78 => wh,
79 => wh,
80 => wh,
81 => wh,
82 => bl,
83 => oa,
84 => bl,
85 => wh,
86 => wh,
87 => wh,
88 => wh,
89 => wh,
90 => wh,
91 => wh,
92 => wh,
93 => wh,
94 => wh,
95 => wh,
96 => wh,
97 => wh,
98 => oa,
99 => bl,
100 => bl,
101 => bl,
102 => wh,
103 => wh,
104 => wh,
105 => wh,
106 => wh,
107 => wh,
108 => wh,
109 => wh,
110 => wh,
111 => wh,
112 => wh,
113 => bu,
114 => wh,
115 => bl,
116 => bl,
117 => bl,
118 => bl,
119 => wh,
120 => bl,
121 => bl,
122 => bl,
123 => bl,
124 => bl,
125 => bl,
126 => wh,
127 => bu,
128 => wh,
129 => bu,
130 => wh,
131 => wh,
132 => bl,
133 => bl,
134 => bl,
135 => bl,
136 => bl,
137 => bl,
138 => bl,
139 => bl,
140 => bl,
141 => bl,
142 => bu,
143 => wh,
144 => bu,
145 => wh,
146 => wh,
147 => wh,
148 => wh,
149 => bl,
150 => bl,
151 => bl,
152 => bl,
153 => bl,
154 => bl,
155 => bl,
156 => bl,
157 => bu,
158 => wh,
159 => wh,
160 => bu,
161 => wh,
162 => wh,
163 => wh,
164 => wh,
165 => wh,
166 => bl,
167 => bl,
168 => bl,
169 => bl,
170 => bl,
171 => bl,
172 => bu,
173 => wh,
174 => wh,
175 => wh,
176 => bu,
177 => wh,
178 => wh,
179 => wh,
180 => wh,
181 => wh,
182 => wh,
183 => bl,
184 => bl,
185 => bl,
186 => wh,
187 => bu,
188 => wh,
189 => wh,
190 => wh,
191 => wh,
192 => bu,
193 => wh,
194 => wh,
195 => wh,
196 => wh,
197 => wh,
198 => wh,
199 => wh,
200 => wh,
201 => wh,
202 => bu,
203 => wh,
204 => wh,
205 => wh,
206 => wh,
207 => wh,
208 => wh,
209 => bu,
210 => wh,
211 => wh,
212 => wh,
213 => wh,
214 => wh,
215 => wh,
216 => wh,
217 => bu,
218 => wh,
219 => wh,
220 => wh,
221 => wh,
222 => wh,
223 => wh,
224 => wh,
225 => wh,
226 => bu,
227 => wh,
228 => wh,
229 => wh,
230 => wh,
231 => bu,
232 => bu,
233 => wh,
234 => wh,
235 => wh,
236 => wh,
237 => wh,
238 => wh,
239 => wh,
240 => wh,
241 => wh,
242 => wh,
243 => bu,
244 => bu,
245 => bu,
246 => bu,
247 => wh,
248 => wh,
249 => wh,
250 => wh,
251 => wh,
252 => wh,
253 => wh,
254 => wh,
255 => wh,
256 => wh,
257 => wh,
258 => wh,
259 => wh,
260 => wh,
261 => wh,
262 => wh,
263 => wh,
264 => wh,
265 => bu,
266 => bu,
267 => bu,
268 => bu,
269 => wh,
270 => wh,
271 => bl,
272 => wh,
273 => wh,
274 => wh,
275 => wh,
276 => wh,
277 => wh,
278 => wh,
279 => bu,
280 => bu,
281 => wh,
282 => wh,
283 => wh,
284 => wh,
285 => bu,
286 => bl,
287 => bl,
288 => wh,
289 => wh,
290 => wh,
291 => wh,
292 => wh,
293 => wh,
294 => bu,
295 => wh,
296 => wh,
297 => wh,
298 => wh,
299 => wh,
300 => wh,
301 => oa,
302 => bl,
303 => bl,
304 => wh,
305 => wh,
306 => wh,
307 => wh,
308 => wh,
309 => bu,
310 => wh,
311 => wh,
312 => wh,
313 => wh,
314 => wh,
315 => wh,
316 => wh,
317 => bl,
318 => oa,
319 => bl,
320 => wh,
321 => wh,
322 => wh,
323 => wh,
324 => bu,
325 => wh,
326 => wh,
327 => wh,
328 => wh,
329 => wh,
330 => wh,
331 => wh,
332 => bl,
333 => bl,
334 => bl,
335 => bu,
336 => wh,
337 => wh,
338 => wh,
339 => bu,
340 => wh,
341 => wh,
342 => wh,
343 => wh,
344 => wh,
345 => wh,
346 => wh,
347 => bl,
348 => bl,
349 => bl,
350 => wh,
351 => bu,
352 => wh,
353 => wh,
354 => bu,
355 => wh,
356 => wh,
357 => wh,
358 => wh,
359 => wh,
360 => wh,
361 => bl,
362 => bl,
363 => bl,
364 => bl,
365 => bl,
366 => wh,
367 => bu,
368 => wh,
369 => bu,
370 => wh,
371 => wh,
372 => wh,
373 => wh,
374 => wh,
375 => bl,
376 => bl,
377 => bl,
378 => bl,
379 => bl,
380 => bl,
381 => wh,
382 => wh,
383 => bu,
384 => bu,
385 => wh,
386 => oa,
387 => oa,
388 => oa,
389 => oa,
390 => bl,
391 => bl,
392 => bl,
393 => bl,
394 => bl,
395 => bl,
396 => wh,
397 => wh,
398 => bu,
399 => wh,
400 => wh,
401 => oa,
402 => bl,
403 => bl,
404 => bl,
405 => bl,
406 => oa,
407 => bl,
408 => bl,
409 => bl,
410 => bl,
411 => wh,
412 => wh,
413 => bu,
414 => wh,
415 => wh,
416 => oa,
417 => bl,
418 => bl,
419 => bl,
420 => bl,
421 => bl,
422 => bl,
423 => oa,
424 => bl,
425 => bl,
426 => bl,
427 => wh,
428 => bu,
429 => wh,
430 => wh,
431 => wh,
432 => oa,
433 => bl,
434 => bl,
435 => bl,
436 => bl,
437 => bl,
438 => bl,
439 => oa,
440 => bl,
441 => bl,
442 => wh,
443 => bu,
444 => wh,
445 => wh,
446 => wh,
447 => wh,
448 => oa,
449 => bl,
450 => bl,
451 => bl,
452 => bl,
453 => bl,
454 => bl,
455 => oa,
456 => bl,
457 => wh,
458 => bu,
459 => wh,
460 => wh,
461 => wh,
462 => wh,
463 => wh,
464 => oa,
465 => bl,
466 => bl,
467 => bl,
468 => bl,
469 => bl,
470 => bl,
471 => oa,
472 => wh,
473 => bu,
474 => wh,
475 => wh,
476 => wh,
477 => wh,
478 => wh,
479 => wh,
480 => bl,
481 => oa,
482 => bl,
483 => bl,
484 => bl,
485 => bl,
486 => oa,
487 => wh,
488 => bu,
489 => wh,
490 => wh,
491 => wh,
492 => wh,
493 => wh,
494 => wh,
495 => wh,
496 => bl,
497 => bl,
498 => oa,
499 => oa,
500 => oa,
501 => oa,
502 => wh,
503 => bu,
504 => wh,
505 => wh,
506 => wh,
507 => wh,
508 => wh,
509 => wh,
510 => wh,
511 => wh,
512 => wh,
513 => wh,
514 => wh,
515 => wh,
516 => wh,
517 => wh,
518 => wh,
519 => bl,
520 => bl,
521 => wh,
522 => wh,
523 => wh,
524 => wh,
525 => wh,
526 => wh,
527 => wh,
528 => wh,
529 => wh,
530 => wh,
531 => wh,
532 => wh,
533 => wh,
534 => wh,
535 => bl,
536 => bl,
537 => bl,
538 => wh,
539 => wh,
540 => wh,
541 => wh,
542 => wh,
543 => wh,
544 => wh,
545 => wh,
546 => wh,
547 => wh,
548 => wh,
549 => wh,
550 => bu,
551 => bl,
552 => bl,
553 => bl,
554 => bu,
555 => wh,
556 => wh,
557 => wh,
558 => bl,
559 => wh,
560 => wh,
561 => wh,
562 => wh,
563 => wh,
564 => wh,
565 => bu,
566 => wh,
567 => wh,
568 => ye,
569 => ye,
570 => wh,
571 => bu,
572 => wh,
573 => wh,
574 => wh,
575 => wh,
576 => wh,
577 => wh,
578 => wh,
579 => wh,
580 => bu,
581 => wh,
582 => wh,
583 => wh,
584 => bl,
585 => bl,
586 => wh,
587 => wh,
588 => bu,
589 => wh,
590 => wh,
591 => wh,
592 => wh,
593 => wh,
594 => wh,
595 => wh,
596 => bu,
597 => wh,
598 => wh,
599 => wh,
600 => bl,
601 => bl,
602 => bl,
603 => wh,
604 => bu,
605 => wh,
606 => wh,
607 => wh,
608 => wh,
609 => wh,
610 => wh,
611 => bu,
612 => wh,
613 => wh,
614 => wh,
615 => wh,
616 => bl,
617 => bl,
618 => bl,
619 => wh,
620 => wh,
621 => bu,
622 => wh,
623 => wh,
624 => wh,
625 => wh,
626 => wh,
627 => bu,
628 => wh,
629 => wh,
630 => wh,
631 => wh,
632 => bl,
633 => bl,
634 => bl,
635 => wh,
636 => wh,
637 => bu,
638 => wh,
639 => wh,
640 => wh,
641 => wh,
642 => wh,
643 => bu,
644 => wh,
645 => wh,
646 => wh,
647 => bl,
648 => bl,
649 => bl,
650 => bl,
651 => wh,
652 => wh,
653 => bu,
654 => wh,
655 => wh,
656 => wh,
657 => wh,
658 => wh,
659 => bu,
660 => wh,
661 => wh,
662 => wh,
663 => bl,
664 => bl,
665 => bl,
666 => bl,
667 => wh,
668 => wh,
669 => bu,
670 => wh,
671 => wh,
672 => wh,
673 => wh,
674 => wh,
675 => bu,
676 => wh,
677 => wh,
678 => bl,
679 => bl,
680 => bl,
681 => bl,
682 => bl,
683 => bl,
684 => wh,
685 => bu,
686 => wh,
687 => wh,
688 => wh,
689 => wh,
690 => wh,
691 => bu,
692 => wh,
693 => wh,
694 => bl,
695 => bl,
696 => bl,
697 => bl,
698 => bl,
699 => bl,
700 => wh,
701 => bu,
702 => wh,
703 => wh,
704 => wh,
705 => wh,
706 => wh,
707 => bu,
708 => wh,
709 => wh,
710 => ye,
711 => ye,
712 => ye,
713 => ye,
714 => bl,
715 => bl,
716 => wh,
717 => bu,
718 => wh,
719 => wh,
720 => wh,
721 => wh,
722 => wh,
723 => bu,
724 => wh,
725 => ye,
726 => bl,
727 => bl,
728 => bl,
729 => bl,
730 => ye,
731 => bl,
732 => wh,
733 => bu,
734 => wh,
735 => wh,
736 => wh,
737 => wh,
738 => wh,
739 => bu,
740 => ye,
741 => bl,
742 => bl,
743 => bl,
744 => bl,
745 => bl,
746 => bl,
747 => ye,
748 => wh,
749 => bu,
750 => wh,
751 => wh,
752 => wh,
753 => wh,
754 => wh,
755 => bu,
756 => ye,
757 => bl,
758 => bl,
759 => bl,
760 => bl,
761 => bl,
762 => bl,
763 => ye,
764 => wh,
765 => bu,
766 => wh,
767 => wh,
768 => wh,
769 => wh,
770 => wh,
771 => bu,
772 => ye,
773 => bl,
774 => bl,
775 => bl,
776 => bl,
777 => bl,
778 => bl,
779 => ye,
780 => wh,
781 => bu,
782 => wh,
783 => wh,
784 => wh,
785 => wh,
786 => wh,
787 => bu,
788 => ye,
789 => bl,
790 => bl,
791 => bl,
792 => bl,
793 => bl,
794 => bl,
795 => ye,
796 => wh,
797 => bu,
798 => wh,
799 => wh,
800 => wh,
801 => wh,
802 => wh,
803 => bu,
804 => wh,
805 => ye,
806 => bl,
807 => bl,
808 => bl,
809 => bl,
810 => ye,
811 => bl,
812 => wh,
813 => bu,
814 => wh,
815 => wh,
816 => wh,
817 => wh,
818 => wh,
819 => bu,
820 => wh,
821 => wh,
822 => ye,
823 => ye,
824 => ye,
825 => ye,
826 => bl,
827 => bl,
828 => wh,
829 => bu,
830 => wh,
831 => wh,
832 => wh,
833 => wh,
834 => wh,
835 => bu,
836 => wh,
837 => wh,
838 => wh,
839 => bl,
840 => bl,
841 => bl,
842 => bl,
843 => bl,
844 => wh,
845 => bu,
846 => wh,
847 => wh,
848 => wh,
849 => wh,
850 => wh,
851 => bu,
852 => wh,
853 => wh,
854 => wh,
855 => bl,
856 => bl,
857 => bl,
858 => bl,
859 => bl,
860 => wh,
861 => bu,
862 => wh,
863 => wh,
864 => wh,
865 => wh,
866 => wh,
867 => bu,
868 => wh,
869 => wh,
870 => wh,
871 => bl,
872 => bl,
873 => bl,
874 => bl,
875 => wh,
876 => wh,
877 => bu,
878 => wh,
879 => wh,
880 => wh,
881 => wh,
882 => wh,
883 => bu,
884 => wh,
885 => wh,
886 => wh,
887 => bl,
888 => bl,
889 => bl,
890 => bl,
891 => wh,
892 => wh,
893 => bu,
894 => wh,
895 => wh,
896 => wh,
897 => wh,
898 => wh,
899 => bu,
900 => wh,
901 => wh,
902 => bl,
903 => bl,
904 => bl,
905 => bl,
906 => wh,
907 => wh,
908 => wh,
909 => bu,
910 => wh,
911 => wh,
912 => wh,
913 => wh,
914 => wh,
915 => bu,
916 => wh,
917 => wh,
918 => bl,
919 => bl,
920 => bl,
921 => bl,
922 => wh,
923 => wh,
924 => wh,
925 => bu,
926 => wh,
927 => wh,
928 => wh,
929 => wh,
930 => wh,
931 => bu,
932 => wh,
933 => bl,
934 => bl,
935 => bl,
936 => bl,
937 => wh,
938 => wh,
939 => wh,
940 => wh,
941 => bu,
942 => wh,
943 => wh,
944 => wh,
945 => wh,
946 => wh,
947 => bu,
948 => bl,
949 => ye,
950 => bl,
951 => bl,
952 => wh,
953 => wh,
954 => wh,
955 => wh,
956 => wh,
957 => bu,
958 => wh,
959 => wh,
960 => wh,
961 => wh,
962 => bl,
963 => bl,
964 => bl,
965 => ye,
966 => bl,
967 => wh,
968 => wh,
969 => wh,
970 => wh,
971 => wh,
972 => bu,
973 => wh,
974 => wh,
975 => wh,
976 => wh,
977 => wh,
978 => bl,
979 => bl,
980 => bl,
981 => wh,
982 => wh,
983 => wh,
984 => wh,
985 => wh,
986 => wh,
987 => wh,
988 => bu,
989 => wh,
990 => wh,
991 => wh,
992 => wh,
993 => wh,
994 => wh,
995 => wh,
996 => wh,
997 => bu,
998 => wh,
999 => wh,
1000 => wh,
1001 => wh,
1002 => wh,
1003 => bu,
1004 => wh,
1005 => wh,
1006 => wh,
1007 => wh,
1008 => wh,
1009 => wh,
1010 => wh,
1011 => wh,
1012 => wh,
1013 => wh,
1014 => bu,
1015 => bu,
1016 => bu,
1017 => bu,
1018 => bu,
1019 => wh,
1020 => wh,
1021 => wh,
1022 => wh,
1023 => wh,
1024 => wh,
1025 => wh,
1026 => wh,
1027 => wh,
1028 => wh,
1029 => wh,
1030 => wh,
1031 => wh,
1032 => wh,
1033 => wh,
1034 => wh,
1035 => wh,
1036 => wh,
1037 => wh,
1038 => wh,
1039 => wh,
1040 => wh,
1041 => wh,
1042 => wh,
1043 => bl,
1044 => bl,
1045 => bl,
1046 => wh,
1047 => wh,
1048 => wh,
1049 => wh,
1050 => wh,
1051 => wh,
1052 => wh,
1053 => wh,
1054 => wh,
1055 => wh,
1056 => wh,
1057 => wh,
1058 => bl,
1059 => wh,
1060 => ye,
1061 => ye,
1062 => bl,
1063 => wh,
1064 => wh,
1065 => wh,
1066 => wh,
1067 => wh,
1068 => wh,
1069 => wh,
1070 => wh,
1071 => wh,
1072 => wh,
1073 => bl,
1074 => lg,
1075 => wh,
1076 => wh,
1077 => lg,
1078 => gr,
1079 => bl,
1080 => bl,
1081 => wh,
1082 => wh,
1083 => wh,
1084 => wh,
1085 => wh,
1086 => wh,
1087 => wh,
1088 => bl,
1089 => wh,
1090 => wh,
1091 => wh,
1092 => wh,
1093 => wh,
1094 => wh,
1095 => wh,
1096 => lg,
1097 => bl,
1098 => wh,
1099 => wh,
1100 => wh,
1101 => wh,
1102 => wh,
1103 => wh,
1104 => bl,
1105 => ge,
1106 => wh,
1107 => ye,
1108 => ye,
1109 => ye,
1110 => ye,
1111 => ye,
1112 => wh,
1113 => ge,
1114 => bl,
1115 => bl,
1116 => wh,
1117 => wh,
1118 => wh,
1119 => wh,
1120 => bl,
1121 => ge,
1122 => wh,
1123 => lg,
1124 => ye,
1125 => oa,
1126 => ye,
1127 => oa,
1128 => wh,
1129 => ge,
1130 => ge,
1131 => ge,
1132 => bl,
1133 => wh,
1134 => wh,
1135 => wh,
1136 => wh,
1137 => bl,
1138 => lg,
1139 => oa,
1140 => ye,
1141 => ye,
1142 => oa,
1143 => ye,
1144 => lg,
1145 => dg,
1146 => dg,
1147 => ge,
1148 => dg,
1149 => bl,
1150 => wh,
1151 => wh,
1152 => wh,
1153 => wh,
1154 => bl,
1155 => oa,
1156 => oa,
1157 => oa,
1158 => lg,
1159 => oa,
1160 => wh,
1161 => wh,
1162 => wh,
1163 => wh,
1164 => wh,
1165 => wh,
1166 => bl,
1167 => wh,
1168 => wh,
1169 => wh,
1170 => wh,
1171 => bl,
1172 => oa,
1173 => oa,
1174 => wh,
1175 => wh,
1176 => wh,
1177 => ge,
1178 => ge,
1179 => ge,
1180 => wh,
1181 => oa,
1182 => oa,
1183 => bl,
1184 => wh,
1185 => wh,
1186 => wh,
1187 => wh,
1188 => bl,
1189 => wh,
1190 => wh,
1191 => wh,
1192 => dg,
1193 => ge,
1194 => dg,
1195 => dg,
1196 => dg,
1197 => wh,
1198 => oa,
1199 => bl,
1200 => wh,
1201 => wh,
1202 => wh,
1203 => wh,
1204 => wh,
1205 => bl,
1206 => wh,
1207 => wh,
1208 => wh,
1209 => wh,
1210 => wh,
1211 => dg,
1212 => dg,
1213 => wh,
1214 => wh,
1215 => bl,
1216 => wh,
1217 => wh,
1218 => wh,
1219 => wh,
1220 => wh,
1221 => wh,
1222 => bl,
1223 => lg,
1224 => gr,
1225 => wh,
1226 => wh,
1227 => dg,
1228 => dg,
1229 => wh,
1230 => bl,
1231 => wh,
1232 => wh,
1233 => wh,
1234 => wh,
1235 => wh,
1236 => wh,
1237 => wh,
1238 => wh,
1239 => bl,
1240 => bl,
1241 => gr,
1242 => ge,
1243 => dg,
1244 => wh,
1245 => lg,
1246 => bl,
1247 => wh,
1248 => wh,
1249 => wh,
1250 => wh,
1251 => wh,
1252 => wh,
1253 => wh,
1254 => wh,
1255 => wh,
1256 => wh,
1257 => bl,
1258 => bl,
1259 => lg,
1260 => wh,
1261 => bl,
1262 => wh,
1263 => wh,
1264 => wh,
1265 => wh,
1266 => wh,
1267 => wh,
1268 => wh,
1269 => wh,
1270 => wh,
1271 => wh,
1272 => wh,
1273 => wh,
1274 => wh,
1275 => bl,
1276 => bl,
1277 => wh,
1278 => wh,
1279 => wh,
1280 => wh,
1281 => wh,
1282 => wh,
1283 => wh,
1284 => wh,
1285 => wh,
1286 => wh,
1287 => wh,
1288 => wh,
1289 => wh,
1290 => wh,
1291 => wh,
1292 => wh,
1293 => wh,
1294 => wh,
1295 => wh,
1296 => wh,
1297 => wh,
1298 => wh,
1299 => wh,
1300 => wh,
1301 => bl,
1302 => bl,
1303 => bl,
1304 => bl,
1305 => bl,
1306 => bl,
1307 => wh,
1308 => wh,
1309 => wh,
1310 => wh,
1311 => wh,
1312 => wh,
1313 => wh,
1314 => wh,
1315 => wh,
1316 => bl,
1317 => ge,
1318 => wh,
1319 => lg,
1320 => wh,
1321 => wh,
1322 => ye,
1323 => bl,
1324 => wh,
1325 => wh,
1326 => wh,
1327 => wh,
1328 => wh,
1329 => wh,
1330 => wh,
1331 => bl,
1332 => ge,
1333 => wh,
1334 => wh,
1335 => ye,
1336 => wh,
1337 => wh,
1338 => lg,
1339 => ye,
1340 => bl,
1341 => wh,
1342 => wh,
1343 => wh,
1344 => wh,
1345 => wh,
1346 => wh,
1347 => bl,
1348 => wh,
1349 => wh,
1350 => wh,
1351 => ye,
1352 => ye,
1353 => wh,
1354 => wh,
1355 => gr,
1356 => bl,
1357 => wh,
1358 => wh,
1359 => wh,
1360 => wh,
1361 => wh,
1362 => wh,
1363 => bl,
1364 => oa,
1365 => oa,
1366 => ye,
1367 => oa,
1368 => ye,
1369 => ye,
1370 => wh,
1371 => lg,
1372 => bl,
1373 => wh,
1374 => wh,
1375 => wh,
1376 => wh,
1377 => wh,
1378 => wh,
1379 => bl,
1380 => oa,
1381 => oa,
1382 => oa,
1383 => ye,
1384 => ye,
1385 => ye,
1386 => wh,
1387 => ge,
1388 => bl,
1389 => wh,
1390 => wh,
1391 => wh,
1392 => wh,
1393 => wh,
1394 => wh,
1395 => bl,
1396 => oa,
1397 => oa,
1398 => ye,
1399 => oa,
1400 => ye,
1401 => wh,
1402 => ge,
1403 => ge,
1404 => bl,
1405 => wh,
1406 => wh,
1407 => wh,
1408 => wh,
1409 => wh,
1410 => wh,
1411 => bl,
1412 => wh,
1413 => wh,
1414 => wh,
1415 => wh,
1416 => wh,
1417 => ge,
1418 => ge,
1419 => ge,
1420 => bl,
1421 => wh,
1422 => wh,
1423 => wh,
1424 => wh,
1425 => wh,
1426 => wh,
1427 => bl,
1428 => wh,
1429 => wh,
1430 => ge,
1431 => ge,
1432 => wh,
1433 => wh,
1434 => dg,
1435 => dg,
1436 => bl,
1437 => wh,
1438 => wh,
1439 => wh,
1440 => wh,
1441 => wh,
1442 => wh,
1443 => bl,
1444 => lg,
1445 => ge,
1446 => wh,
1447 => ge,
1448 => ge,
1449 => wh,
1450 => wh,
1451 => dg,
1452 => bl,
1453 => wh,
1454 => wh,
1455 => wh,
1456 => wh,
1457 => wh,
1458 => wh,
1459 => bl,
1460 => gr,
1461 => wh,
1462 => wh,
1463 => dg,
1464 => ge,
1465 => wh,
1466 => wh,
1467 => wh,
1468 => bl,
1469 => wh,
1470 => wh,
1471 => wh,
1472 => wh,
1473 => wh,
1474 => wh,
1475 => bl,
1476 => lg,
1477 => dg,
1478 => dg,
1479 => dg,
1480 => dg,
1481 => wh,
1482 => oa,
1483 => oa,
1484 => bl,
1485 => wh,
1486 => wh,
1487 => wh,
1488 => wh,
1489 => wh,
1490 => wh,
1491 => wh,
1492 => bl,
1493 => lg,
1494 => dg,
1495 => dg,
1496 => lg,
1497 => wh,
1498 => oa,
1499 => bl,
1500 => wh,
1501 => wh,
1502 => wh,
1503 => wh,
1504 => wh,
1505 => wh,
1506 => wh,
1507 => wh,
1508 => wh,
1509 => bl,
1510 => bl,
1511 => bl,
1512 => bl,
1513 => bl,
1514 => bl,
1515 => wh,
1516 => wh,
1517 => wh,
1518 => wh,
1519 => wh,
1520 => wh,
1521 => wh,
1522 => wh,
1523 => wh,
1524 => wh,
1525 => wh,
1526 => wh,
1527 => wh,
1528 => wh,
1529 => wh,
1530 => wh,
1531 => wh,
1532 => wh,
1533 => wh,
1534 => wh,
1535 => wh,
1536 => wh,
1537 => wh,
1538 => wh,
1539 => wh,
1540 => wh,
1541 => wh,
1542 => wh,
1543 => wh,
1544 => wh,
1545 => wh,
1546 => wh,
1547 => wh,
1548 => wh,
1549 => wh,
1550 => wh,
1551 => wh,
1552 => wh,
1553 => wh,
1554 => wh,
1555 => wh,
1556 => wh,
1557 => wh,
1558 => wh,
1559 => wh,
1560 => wh,
1561 => wh,
1562 => wh,
1563 => bl,
1564 => bl,
1565 => wh,
1566 => wh,
1567 => wh,
1568 => wh,
1569 => wh,
1570 => wh,
1571 => wh,
1572 => wh,
1573 => wh,
1574 => wh,
1575 => wh,
1576 => wh,
1577 => wh,
1578 => bl,
1579 => ge,
1580 => ge,
1581 => bl,
1582 => wh,
1583 => wh,
1584 => wh,
1585 => wh,
1586 => wh,
1587 => wh,
1588 => wh,
1589 => wh,
1590 => wh,
1591 => wh,
1592 => bl,
1593 => bl,
1594 => wh,
1595 => wh,
1596 => wh,
1597 => wh,
1598 => bl,
1599 => wh,
1600 => wh,
1601 => wh,
1602 => wh,
1603 => wh,
1604 => wh,
1605 => wh,
1606 => bl,
1607 => bl,
1608 => oa,
1609 => oa,
1610 => oa,
1611 => ye,
1612 => ye,
1613 => wh,
1614 => lg,
1615 => bl,
1616 => wh,
1617 => wh,
1618 => wh,
1619 => wh,
1620 => wh,
1621 => bl,
1622 => wh,
1623 => oa,
1624 => oa,
1625 => ye,
1626 => ye,
1627 => ye,
1628 => ye,
1629 => wh,
1630 => wh,
1631 => bl,
1632 => wh,
1633 => wh,
1634 => wh,
1635 => bl,
1636 => bl,
1637 => wh,
1638 => wh,
1639 => wh,
1640 => oa,
1641 => oa,
1642 => oa,
1643 => ye,
1644 => ye,
1645 => wh,
1646 => ye,
1647 => bl,
1648 => wh,
1649 => wh,
1650 => bl,
1651 => wh,
1652 => lg,
1653 => ge,
1654 => wh,
1655 => wh,
1656 => lg,
1657 => oa,
1658 => ye,
1659 => ye,
1660 => wh,
1661 => lg,
1662 => ye,
1663 => bl,
1664 => wh,
1665 => bl,
1666 => gr,
1667 => lg,
1668 => wh,
1669 => dg,
1670 => ge,
1671 => wh,
1672 => oa,
1673 => ye,
1674 => oa,
1675 => ye,
1676 => wh,
1677 => gr,
1678 => bl,
1679 => wh,
1680 => bl,
1681 => lg,
1682 => dg,
1683 => wh,
1684 => wh,
1685 => ge,
1686 => dg,
1687 => wh,
1688 => wh,
1689 => wh,
1690 => wh,
1691 => wh,
1692 => wh,
1693 => bl,
1694 => wh,
1695 => wh,
1696 => bl,
1697 => lg,
1698 => dg,
1699 => ge,
1700 => ge,
1701 => dg,
1702 => ge,
1703 => wh,
1704 => dg,
1705 => ge,
1706 => ge,
1707 => lg,
1708 => bl,
1709 => wh,
1710 => wh,
1711 => wh,
1712 => bl,
1713 => wh,
1714 => wh,
1715 => dg,
1716 => dg,
1717 => ge,
1718 => wh,
1719 => wh,
1720 => ge,
1721 => dg,
1722 => bl,
1723 => bl,
1724 => wh,
1725 => wh,
1726 => wh,
1727 => wh,
1728 => wh,
1729 => bl,
1730 => lg,
1731 => wh,
1732 => wh,
1733 => wh,
1734 => wh,
1735 => wh,
1736 => dg,
1737 => bl,
1738 => wh,
1739 => wh,
1740 => wh,
1741 => wh,
1742 => wh,
1743 => wh,
1744 => wh,
1745 => wh,
1746 => bl,
1747 => wh,
1748 => wh,
1749 => oa,
1750 => wh,
1751 => dg,
1752 => bl,
1753 => wh,
1754 => wh,
1755 => wh,
1756 => wh,
1757 => wh,
1758 => wh,
1759 => wh,
1760 => wh,
1761 => wh,
1762 => wh,
1763 => bl,
1764 => oa,
1765 => oa,
1766 => bl,
1767 => bl,
1768 => wh,
1769 => wh,
1770 => wh,
1771 => wh,
1772 => wh,
1773 => wh,
1774 => wh,
1775 => wh,
1776 => wh,
1777 => wh,
1778 => wh,
1779 => wh,
1780 => bl,
1781 => bl,
1782 => wh,
1783 => wh,
1784 => wh,
1785 => wh,
1786 => wh,
1787 => wh,
1788 => wh,
1789 => wh,
1790 => wh,
1791 => wh,
1792 => wh,
1793 => wh,
1794 => wh,
1795 => wh,
1796 => wh,
1797 => wh,
1798 => wh,
1799 => wh,
1800 => wh,
1801 => wh,
1802 => wh,
1803 => wh,
1804 => wh,
1805 => wh,
1806 => wh,
1807 => wh,
1808 => wh,
1809 => wh,
1810 => wh,
1811 => wh,
1812 => wh,
1813 => wh,
1814 => wh,
1815 => wh,
1816 => wh,
1817 => wh,
1818 => wh,
1819 => wh,
1820 => wh,
1821 => wh,
1822 => wh,
1823 => wh,
1824 => wh,
1825 => wh,
1826 => wh,
1827 => wh,
1828 => wh,
1829 => wh,
1830 => wh,
1831 => wh,
1832 => wh,
1833 => wh,
1834 => wh,
1835 => wh,
1836 => wh,
1837 => wh,
1838 => wh,
1839 => wh,
1840 => wh,
1841 => wh,
1842 => bl,
1843 => bl,
1844 => bl,
1845 => bl,
1846 => bl,
1847 => bl,
1848 => bl,
1849 => bl,
1850 => bl,
1851 => bl,
1852 => bl,
1853 => bl,
1854 => wh,
1855 => wh,
1856 => wh,
1857 => bl,
1858 => ye,
1859 => lg,
1860 => gr,
1861 => wh,
1862 => ge,
1863 => ge,
1864 => dg,
1865 => ge,
1866 => dg,
1867 => wh,
1868 => wh,
1869 => oa,
1870 => bl,
1871 => wh,
1872 => bl,
1873 => ye,
1874 => wh,
1875 => lg,
1876 => wh,
1877 => ye,
1878 => wh,
1879 => ge,
1880 => dg,
1881 => dg,
1882 => wh,
1883 => wh,
1884 => wh,
1885 => oa,
1886 => oa,
1887 => bl,
1888 => bl,
1889 => wh,
1890 => wh,
1891 => wh,
1892 => ye,
1893 => ye,
1894 => ye,
1895 => wh,
1896 => ge,
1897 => wh,
1898 => wh,
1899 => wh,
1900 => wh,
1901 => wh,
1902 => wh,
1903 => bl,
1904 => bl,
1905 => lg,
1906 => wh,
1907 => ye,
1908 => ye,
1909 => oa,
1910 => oa,
1911 => ye,
1912 => wh,
1913 => wh,
1914 => ge,
1915 => ge,
1916 => dg,
1917 => dg,
1918 => wh,
1919 => bl,
1920 => bl,
1921 => wh,
1922 => ye,
1923 => ye,
1924 => oa,
1925 => ye,
1926 => oa,
1927 => ye,
1928 => wh,
1929 => ge,
1930 => dg,
1931 => dg,
1932 => ge,
1933 => dg,
1934 => lg,
1935 => bl,
1936 => bl,
1937 => ge,
1938 => wh,
1939 => wh,
1940 => ye,
1941 => oa,
1942 => oa,
1943 => wh,
1944 => wh,
1945 => ge,
1946 => dg,
1947 => wh,
1948 => wh,
1949 => dg,
1950 => dg,
1951 => bl,
1952 => bl,
1953 => ge,
1954 => wh,
1955 => wh,
1956 => oa,
1957 => oa,
1958 => oa,
1959 => wh,
1960 => wh,
1961 => ge,
1962 => dg,
1963 => wh,
1964 => wh,
1965 => dg,
1966 => dg,
1967 => bl,
1968 => wh,
1969 => bl,
1970 => dg,
1971 => wh,
1972 => oa,
1973 => oa,
1974 => oa,
1975 => wh,
1976 => wh,
1977 => wh,
1978 => dg,
1979 => lg,
1980 => gr,
1981 => lg,
1982 => bl,
1983 => wh,
1984 => wh,
1985 => wh,
1986 => bl,
1987 => bl,
1988 => bl,
1989 => bl,
1990 => bl,
1991 => bl,
1992 => bl,
1993 => bl,
1994 => bl,
1995 => bl,
1996 => bl,
1997 => bl,
1998 => wh,
1999 => wh,
2000 => wh,
2001 => wh,
2002 => wh,
2003 => wh,
2004 => wh,
2005 => wh,
2006 => wh,
2007 => wh,
2008 => wh,
2009 => wh,
2010 => wh,
2011 => wh,
2012 => wh,
2013 => wh,
2014 => wh,
2015 => wh,
2016 => wh,
2017 => wh,
2018 => wh,
2019 => wh,
2020 => wh,
2021 => wh,
2022 => wh,
2023 => wh,
2024 => wh,
2025 => wh,
2026 => wh,
2027 => wh,
2028 => wh,
2029 => wh,
2030 => wh,
2031 => wh,
2032 => wh,
2033 => wh,
2034 => wh,
2035 => wh,
2036 => wh,
2037 => wh,
2038 => wh,
2039 => wh,
2040 => wh,
2041 => wh,
2042 => wh,
2043 => wh,
2044 => wh,
2045 => wh,
2046 => wh,
2047 => wh
    ); 
    
    attribute ram_style : string;
    attribute ram_style of tile_data_map_d : signal is "block";
begin
    
      process(i_tile_id, i_x, i_y)
          variable readIndex : std_logic_vector (10 downto 0);
          variable readIndex_int : integer;
          begin
          readIndex := i_tile_id & i_y & i_x;
          readIndex_int := to_integer(unsigned(readIndex));
          o_colorCode <= tile_data_map_d(readIndex_int);
      end process;
      
      process(i_clk)
      variable writeIndex : std_logic_vector (10 downto 0);
      variable writeIndex_int : integer;
      begin
        if rising_edge(i_clk) then
            if i_ch_we = '1' then
                writeIndex := i_tile_id_write & i_ch_y & i_ch_x;
                writeIndex_int := to_integer(unsigned(writeIndex));
                tile_data_map_d(writeIndex_int) <= i_ch_cc;
            end if;
        end if;
      end process;

end Behavioral;
