library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity TuileBackBuff2 is
    Port(
    i_x : in STD_LOGIC_VECTOR (2 downto 0);
    i_y : in STD_LOGIC_VECTOR (2 downto 0);
    i_tile_id : in STD_LOGIC_VECTOR (4 downto 0);
    i_ch_x : in STD_LOGIC_VECTOR (2 downto 0);
    i_ch_y : in STD_LOGIC_VECTOR (2 downto 0);
    i_ch_cc : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_we : in std_logic;
    i_clk : in STD_LOGIC;
    i_flip_y : in STD_LOGIC;
    i_tile_id_write : in STD_LOGIC_VECTOR (4 downto 0);
    o_colorCode : out STD_LOGIC_VECTOR (3 downto 0));
end TuileBackBuff2;

architecture Behavioral of TuileBackBuff2 is
constant wh : std_logic_vector (3 downto 0) := "0000"; -- White
constant bl : std_logic_vector (3 downto 0) := "0001"; -- Black
constant ye : std_logic_vector (3 downto 0) := "0010"; -- Yellow
constant dg : std_logic_vector (3 downto 0) := "0011"; -- Dark Green
constant oa : std_logic_vector (3 downto 0) := "0100"; -- Orange
constant bu : std_logic_vector (3 downto 0) := "0101"; -- Blue
constant ge : std_logic_vector (3 downto 0) := "0110"; -- Green
constant lo : std_logic_vector (3 downto 0) := "0111"; -- Light Brown
constant br : std_logic_vector (3 downto 0) := "1000"; -- Brown
constant lg : std_logic_vector (3 downto 0) := "1001"; -- Light Gray
constant gr : std_logic_vector (3 downto 0) := "1010"; -- Gray
constant lb : std_logic_vector (3 downto 0) := "1011"; -- Light Blue
constant sb : std_logic_vector (3 downto 0) := "1100"; -- Sky Blue
constant sa : std_logic_vector (3 downto 0) := "1101"; -- Salmon
constant pi : std_logic_vector (3 downto 0) := "1110"; -- Pink
constant pu : std_logic_vector (3 downto 0) := "1111"; -- Purple

    type tuile_out_array_t is array (0 to 31) of std_logic_vector(3 downto 0);
    signal tuile_outputs : tuile_out_array_t;
    signal tuile_write_enable : std_logic_vector(31 downto 0);
    
    type tile_d_array_t is array (0 to 1023) of std_logic_vector(3 downto 0);
    signal tile_data_map_d : tile_d_array_t :=
    (
        0 => wh,
        1 => wh,
        2 => wh,
        3 => wh,
        4 => wh,
        5 => wh,
        6 => wh,
        7 => wh,
        8 => wh,
        9 => wh,
        10 => wh,
        11 => wh,
        12 => wh,
        13 => wh,
        14 => wh,
        15 => wh,
        16 => wh,
        17 => wh,
        18 => wh,
        19 => wh,
        20 => wh,
        21 => wh,
        22 => wh,
        23 => wh,
        24 => wh,
        25 => wh,
        26 => wh,
        27 => wh,
        28 => wh,
        29 => wh,
        30 => wh,
        31 => wh,
        32 => wh,
        33 => wh,
        34 => wh,
        35 => wh,
        36 => wh,
        37 => wh,
        38 => wh,
        39 => wh,
        40 => wh,
        41 => wh,
        42 => wh,
        43 => wh,
        44 => wh,
        45 => wh,
        46 => wh,
        47 => wh,
        48 => wh,
        49 => wh,
        50 => wh,
        51 => wh,
        52 => wh,
        53 => wh,
        54 => wh,
        55 => wh,
        56 => wh,
        57 => wh,
        58 => wh,
        59 => wh,
        60 => wh,
        61 => wh,
        62 => wh,
        63 => wh,
        64 => wh,
        65 => wh,
        66 => sb,
        67 => lb,
        68 => lb,
        69 => sb,
        70 => wh,
        71 => wh,
        72 => wh,
        73 => wh,
        74 => sb,
        75 => lb,
        76 => lb,
        77 => sb,
        78 => sb,
        79 => wh,
        80 => wh,
        81 => wh,
        82 => sb,
        83 => lb,
        84 => lb,
        85 => sb,
        86 => wh,
        87 => wh,
        88 => wh,
        89 => sb,
        90 => lb,
        91 => lb,
        92 => lb,
        93 => sb,
        94 => wh,
        95 => wh,
        96 => wh,
        97 => wh,
        98 => sb,
        99 => lb,
        100 => lb,
        101 => sb,
        102 => wh,
        103 => wh,
        104 => wh,
        105 => wh,
        106 => sb,
        107 => lb,
        108 => lb,
        109 => sb,
        110 => sb,
        111 => wh,
        112 => wh,
        113 => sb,
        114 => sb,
        115 => lb,
        116 => lb,
        117 => sb,
        118 => wh,
        119 => wh,
        120 => wh,
        121 => wh,
        122 => sb,
        123 => lb,
        124 => lb,
        125 => sb,
        126 => wh,
        127 => wh,
        128 => wh,
        129 => wh,
        130 => pi,
        131 => sa,
        132 => sa,
        133 => pi,
        134 => wh,
        135 => wh,
        136 => wh,
        137 => wh,
        138 => pi,
        139 => sa,
        140 => sa,
        141 => pi,
        142 => wh,
        143 => wh,
        144 => wh,
        145 => pi,
        146 => pi,
        147 => sa,
        148 => sa,
        149 => pi,
        150 => wh,
        151 => wh,
        152 => wh,
        153 => wh,
        154 => pi,
        155 => sa,
        156 => sa,
        157 => pi,
        158 => wh,
        159 => wh,
        160 => wh,
        161 => wh,
        162 => pi,
        163 => sa,
        164 => sa,
        165 => sa,
        166 => pi,
        167 => wh,
        168 => wh,
        169 => wh,
        170 => pi,
        171 => sa,
        172 => sa,
        173 => pi,
        174 => wh,
        175 => wh,
        176 => wh,
        177 => pi,
        178 => pi,
        179 => sa,
        180 => sa,
        181 => pi,
        182 => wh,
        183 => wh,
        184 => wh,
        185 => wh,
        186 => pi,
        187 => sa,
        188 => sa,
        189 => pi,
        190 => wh,
        191 => wh,
        192 => wh,
        193 => wh,
        194 => wh,
        195 => wh,
        196 => wh,
        197 => wh,
        198 => wh,
        199 => wh,
        200 => wh,
        201 => wh,
        202 => wh,
        203 => wh,
        204 => wh,
        205 => lg,
        206 => lg,
        207 => pi,
        208 => wh,
        209 => wh,
        210 => wh,
        211 => lg,
        212 => lg,
        213 => lg,
        214 => lg,
        215 => wh,
        216 => wh,
        217 => wh,
        218 => lg,
        219 => lg,
        220 => lg,
        221 => wh,
        222 => gr,
        223 => lg,
        224 => wh,
        225 => wh,
        226 => lg,
        227 => lg,
        228 => gr,
        229 => lg,
        230 => lg,
        231 => lg,
        232 => wh,
        233 => lg,
        234 => wh,
        235 => gr,
        236 => wh,
        237 => gr,
        238 => lg,
        239 => lg,
        240 => wh,
        241 => wh,
        242 => wh,
        243 => wh,
        244 => lg,
        245 => gr,
        246 => lg,
        247 => wh,
        248 => wh,
        249 => wh,
        250 => wh,
        251 => wh,
        252 => wh,
        253 => wh,
        254 => wh,
        255 => lg,
        256 => lg,
        257 => lg,
        258 => wh,
        259 => lg,
        260 => lg,
        261 => lg,
        262 => lg,
        263 => wh,
        264 => wh,
        265 => wh,
        266 => wh,
        267 => pi,
        268 => wh,
        269 => pi,
        270 => wh,
        271 => lg,
        272 => wh,
        273 => pi,
        274 => wh,
        275 => pi,
        276 => pi,
        277 => wh,
        278 => pi,
        279 => pi,
        280 => lg,
        281 => wh,
        282 => lg,
        283 => pi,
        284 => gr,
        285 => pi,
        286 => lg,
        287 => gr,
        288 => pi,
        289 => lg,
        290 => lg,
        291 => gr,
        292 => gr,
        293 => gr,
        294 => gr,
        295 => lg,
        296 => gr,
        297 => gr,
        298 => gr,
        299 => lg,
        300 => gr,
        301 => gr,
        302 => lg,
        303 => gr,
        304 => wh,
        305 => gr,
        306 => gr,
        307 => gr,
        308 => pi,
        309 => gr,
        310 => gr,
        311 => gr,
        312 => wh,
        313 => wh,
        314 => wh,
        315 => wh,
        316 => gr,
        317 => wh,
        318 => gr,
        319 => pi,
        320 => wh,
        321 => wh,
        322 => wh,
        323 => wh,
        324 => wh,
        325 => wh,
        326 => wh,
        327 => wh,
        328 => lg,
        329 => lg,
        330 => wh,
        331 => wh,
        332 => wh,
        333 => wh,
        334 => wh,
        335 => wh,
        336 => gr,
        337 => gr,
        338 => gr,
        339 => gr,
        340 => wh,
        341 => wh,
        342 => wh,
        343 => wh,
        344 => pi,
        345 => pi,
        346 => lg,
        347 => gr,
        348 => gr,
        349 => wh,
        350 => wh,
        351 => wh,
        352 => pi,
        353 => gr,
        354 => gr,
        355 => lg,
        356 => lg,
        357 => wh,
        358 => wh,
        359 => wh,
        360 => gr,
        361 => lg,
        362 => gr,
        363 => gr,
        364 => lg,
        365 => gr,
        366 => wh,
        367 => wh,
        368 => gr,
        369 => gr,
        370 => pi,
        371 => lg,
        372 => pi,
        373 => gr,
        374 => wh,
        375 => wh,
        376 => gr,
        377 => pi,
        378 => pi,
        379 => wh,
        380 => wh,
        381 => pi,
        382 => wh,
        383 => wh,
        384 => wh,
        385 => wh,
        386 => wh,
        387 => wh,
        388 => wh,
        389 => wh,
        390 => wh,
        391 => wh,
        392 => wh,
        393 => wh,
        394 => wh,
        395 => pi,
        396 => lg,
        397 => pi,
        398 => lg,
        399 => wh,
        400 => wh,
        401 => wh,
        402 => pi,
        403 => wh,
        404 => lg,
        405 => pi,
        406 => wh,
        407 => pi,
        408 => wh,
        409 => pi,
        410 => lg,
        411 => pi,
        412 => lg,
        413 => lg,
        414 => lg,
        415 => wh,
        416 => wh,
        417 => lg,
        418 => wh,
        419 => lg,
        420 => lg,
        421 => lg,
        422 => lg,
        423 => lg,
        424 => lg,
        425 => lg,
        426 => lg,
        427 => pi,
        428 => lg,
        429 => lg,
        430 => wh,
        431 => lg,
        432 => wh,
        433 => lg,
        434 => pi,
        435 => lg,
        436 => gr,
        437 => pi,
        438 => lg,
        439 => gr,
        440 => lg,
        441 => lg,
        442 => lg,
        443 => lg,
        444 => lg,
        445 => lg,
        446 => gr,
        447 => gr,
        448 => lg,
        449 => wh,
        450 => lg,
        451 => lg,
        452 => pi,
        453 => gr,
        454 => gr,
        455 => gr,
        456 => wh,
        457 => pi,
        458 => gr,
        459 => lg,
        460 => gr,
        461 => lg,
        462 => gr,
        463 => gr,
        464 => lg,
        465 => lg,
        466 => lg,
        467 => gr,
        468 => gr,
        469 => gr,
        470 => lg,
        471 => pi,
        472 => lg,
        473 => gr,
        474 => gr,
        475 => gr,
        476 => gr,
        477 => lg,
        478 => gr,
        479 => lg,
        480 => lg,
        481 => pi,
        482 => gr,
        483 => gr,
        484 => gr,
        485 => gr,
        486 => lg,
        487 => gr,
        488 => lg,
        489 => pi,
        490 => gr,
        491 => gr,
        492 => lg,
        493 => lg,
        494 => gr,
        495 => lg,
        496 => wh,
        497 => gr,
        498 => wh,
        499 => lg,
        500 => gr,
        501 => pi,
        502 => gr,
        503 => pi,
        504 => wh,
        505 => wh,
        506 => gr,
        507 => wh,
        508 => wh,
        509 => gr,
        510 => wh,
        511 => wh,
        512 => pi,
        513 => wh,
        514 => pi,
        515 => pi,
        516 => pi,
        517 => gr,
        518 => wh,
        519 => wh,
        520 => lg,
        521 => gr,
        522 => pi,
        523 => lg,
        524 => gr,
        525 => gr,
        526 => gr,
        527 => wh,
        528 => gr,
        529 => gr,
        530 => gr,
        531 => gr,
        532 => gr,
        533 => gr,
        534 => gr,
        535 => gr,
        536 => lg,
        537 => gr,
        538 => lg,
        539 => gr,
        540 => gr,
        541 => gr,
        542 => gr,
        543 => wh,
        544 => lg,
        545 => gr,
        546 => gr,
        547 => gr,
        548 => lg,
        549 => gr,
        550 => wh,
        551 => gr,
        552 => gr,
        553 => gr,
        554 => gr,
        555 => gr,
        556 => gr,
        557 => gr,
        558 => gr,
        559 => wh,
        560 => wh,
        561 => gr,
        562 => lg,
        563 => gr,
        564 => pi,
        565 => pi,
        566 => pi,
        567 => gr,
        568 => wh,
        569 => pi,
        570 => wh,
        571 => pi,
        572 => pi,
        573 => wh,
        574 => wh,
        575 => pi,
        576 => wh,
        577 => wh,
        578 => sb,
        579 => lb,
        580 => lb,
        581 => sb,
        582 => wh,
        583 => wh,
        584 => wh,
        585 => wh,
        586 => sb,
        587 => sb,
        588 => lb,
        589 => sb,
        590 => wh,
        591 => wh,
        592 => wh,
        593 => wh,
        594 => wh,
        595 => lb,
        596 => lb,
        597 => wh,
        598 => wh,
        599 => wh,
        600 => wh,
        601 => wh,
        602 => wh,
        603 => sb,
        604 => lb,
        605 => wh,
        606 => wh,
        607 => wh,
        608 => wh,
        609 => wh,
        610 => sb,
        611 => wh,
        612 => sb,
        613 => wh,
        614 => wh,
        615 => wh,
        616 => wh,
        617 => wh,
        618 => wh,
        619 => lb,
        620 => sb,
        621 => wh,
        622 => wh,
        623 => wh,
        624 => wh,
        625 => wh,
        626 => wh,
        627 => sb,
        628 => wh,
        629 => wh,
        630 => wh,
        631 => wh,
        632 => wh,
        633 => wh,
        634 => wh,
        635 => wh,
        636 => wh,
        637 => wh,
        638 => wh,
        639 => wh,
        640 => wh,
        641 => wh,
        642 => pi,
        643 => sa,
        644 => pi,
        645 => pi,
        646 => wh,
        647 => wh,
        648 => wh,
        649 => wh,
        650 => pi,
        651 => sa,
        652 => sa,
        653 => pi,
        654 => wh,
        655 => wh,
        656 => wh,
        657 => wh,
        658 => pi,
        659 => pi,
        660 => sa,
        661 => pi,
        662 => wh,
        663 => wh,
        664 => wh,
        665 => wh,
        666 => wh,
        667 => sa,
        668 => pi,
        669 => wh,
        670 => wh,
        671 => wh,
        672 => wh,
        673 => wh,
        674 => wh,
        675 => pi,
        676 => pi,
        677 => wh,
        678 => wh,
        679 => wh,
        680 => wh,
        681 => wh,
        682 => wh,
        683 => wh,
        684 => sa,
        685 => wh,
        686 => wh,
        687 => wh,
        688 => wh,
        689 => wh,
        690 => wh,
        691 => wh,
        692 => wh,
        693 => wh,
        694 => wh,
        695 => wh,
        696 => wh,
        697 => wh,
        698 => wh,
        699 => pi,
        700 => wh,
        701 => wh,
        702 => wh,
        703 => wh,
        704 => bl,
        705 => bl,
        706 => bl,
        707 => bl,
        708 => bl,
        709 => bl,
        710 => bl,
        711 => bl,
        712 => bl,
        713 => bl,
        714 => bl,
        715 => bl,
        716 => bl,
        717 => bl,
        718 => bl,
        719 => bl,
        720 => bl,
        721 => bl,
        722 => bl,
        723 => bl,
        724 => bl,
        725 => bl,
        726 => bl,
        727 => bl,
        728 => bl,
        729 => bl,
        730 => bl,
        731 => bl,
        732 => bl,
        733 => bl,
        734 => bl,
        735 => bl,
        736 => bl,
        737 => bl,
        738 => bl,
        739 => bl,
        740 => bl,
        741 => bl,
        742 => bl,
        743 => bl,
        744 => bl,
        745 => bl,
        746 => bl,
        747 => bl,
        748 => bl,
        749 => bl,
        750 => bl,
        751 => bl,
        752 => bl,
        753 => bl,
        754 => bl,
        755 => bl,
        756 => bl,
        757 => bl,
        758 => bl,
        759 => bl,
        760 => bl,
        761 => bl,
        762 => bl,
        763 => bl,
        764 => bl,
        765 => bl,
        766 => bl,
        767 => bl,
        768 => ye,
        769 => ye,
        770 => ye,
        771 => ye,
        772 => dg,
        773 => dg,
        774 => dg,
        775 => dg,
        776 => ye,
        777 => ye,
        778 => ye,
        779 => ye,
        780 => dg,
        781 => dg,
        782 => dg,
        783 => dg,
        784 => ye,
        785 => ye,
        786 => ye,
        787 => ye,
        788 => dg,
        789 => dg,
        790 => dg,
        791 => dg,
        792 => ye,
        793 => ye,
        794 => ye,
        795 => ye,
        796 => dg,
        797 => dg,
        798 => dg,
        799 => dg,
        800 => ye,
        801 => ye,
        802 => ye,
        803 => ye,
        804 => dg,
        805 => dg,
        806 => dg,
        807 => dg,
        808 => ye,
        809 => ye,
        810 => ye,
        811 => ye,
        812 => dg,
        813 => dg,
        814 => dg,
        815 => dg,
        816 => ye,
        817 => ye,
        818 => ye,
        819 => ye,
        820 => dg,
        821 => dg,
        822 => dg,
        823 => dg,
        824 => ye,
        825 => ye,
        826 => ye,
        827 => ye,
        828 => dg,
        829 => dg,
        830 => dg,
        831 => dg,
        832 => oa,
        833 => oa,
        834 => oa,
        835 => oa,
        836 => bu,
        837 => bu,
        838 => bu,
        839 => bu,
        840 => oa,
        841 => oa,
        842 => oa,
        843 => oa,
        844 => bu,
        845 => bu,
        846 => bu,
        847 => bu,
        848 => oa,
        849 => oa,
        850 => oa,
        851 => oa,
        852 => bu,
        853 => bu,
        854 => bu,
        855 => bu,
        856 => oa,
        857 => oa,
        858 => oa,
        859 => oa,
        860 => bu,
        861 => bu,
        862 => bu,
        863 => bu,
        864 => oa,
        865 => oa,
        866 => oa,
        867 => oa,
        868 => bu,
        869 => bu,
        870 => bu,
        871 => bu,
        872 => oa,
        873 => oa,
        874 => oa,
        875 => oa,
        876 => bu,
        877 => bu,
        878 => bu,
        879 => bu,
        880 => oa,
        881 => oa,
        882 => oa,
        883 => oa,
        884 => bu,
        885 => bu,
        886 => bu,
        887 => bu,
        888 => oa,
        889 => oa,
        890 => oa,
        891 => oa,
        892 => bu,
        893 => bu,
        894 => bu,
        895 => bu,
        896 => ge,
        897 => ge,
        898 => ge,
        899 => ge,
        900 => pu,
        901 => pu,
        902 => pu,
        903 => pu,
        904 => ge,
        905 => ge,
        906 => ge,
        907 => ge,
        908 => pu,
        909 => pu,
        910 => pu,
        911 => pu,
        912 => ge,
        913 => ge,
        914 => ge,
        915 => ge,
        916 => pu,
        917 => pu,
        918 => pu,
        919 => pu,
        920 => ge,
        921 => ge,
        922 => ge,
        923 => ge,
        924 => pu,
        925 => pu,
        926 => pu,
        927 => pu,
        928 => ge,
        929 => ge,
        930 => ge,
        931 => ge,
        932 => pu,
        933 => pu,
        934 => pu,
        935 => pu,
        936 => ge,
        937 => ge,
        938 => ge,
        939 => ge,
        940 => pu,
        941 => pu,
        942 => pu,
        943 => pu,
        944 => ge,
        945 => ge,
        946 => ge,
        947 => ge,
        948 => pu,
        949 => pu,
        950 => pu,
        951 => pu,
        952 => ge,
        953 => ge,
        954 => ge,
        955 => ge,
        956 => pu,
        957 => pu,
        958 => pu,
        959 => pu,
        960 => lo,
        961 => lo,
        962 => lo,
        963 => lo,
        964 => br,
        965 => br,
        966 => br,
        967 => br,
        968 => lo,
        969 => lo,
        970 => lo,
        971 => lo,
        972 => br,
        973 => br,
        974 => br,
        975 => br,
        976 => lo,
        977 => lo,
        978 => lo,
        979 => lo,
        980 => br,
        981 => br,
        982 => br,
        983 => br,
        984 => lo,
        985 => lo,
        986 => lo,
        987 => lo,
        988 => br,
        989 => br,
        990 => br,
        991 => br,
        992 => lo,
        993 => lo,
        994 => lo,
        995 => lo,
        996 => br,
        997 => br,
        998 => br,
        999 => br,
        1000 => lo,
        1001 => lo,
        1002 => lo,
        1003 => lo,
        1004 => br,
        1005 => br,
        1006 => br,
        1007 => br,
        1008 => lo,
        1009 => lo,
        1010 => lo,
        1011 => lo,
        1012 => br,
        1013 => br,
        1014 => br,
        1015 => br,
        1016 => lo,
        1017 => lo,
        1018 => lo,
        1019 => lo,
        1020 => br,
        1021 => br,
        1022 => br,
        1023 => br
    ); 
    
    attribute ram_style : string;
    attribute ram_style of tile_data_map_d : signal is "block";
begin
    
      process(i_tile_id, i_x, i_y)
          variable readIndex : std_logic_vector (10 downto 0);
          variable readIndex_int : integer;
          begin
          readIndex := i_tile_id & i_y & i_x;
          readIndex_int := to_integer(unsigned(readIndex));
          o_colorCode <= tile_data_map_d(readIndex_int);
      end process;
      
      process(i_clk)
      variable writeIndex : std_logic_vector (10 downto 0);
      variable writeIndex_int : integer;
      begin
        if rising_edge(i_clk) then
            if i_ch_we = '1' then
                writeIndex := i_tile_id_write & i_ch_y & i_ch_x;
                writeIndex_int := to_integer(unsigned(writeIndex));
                tile_data_map_d(writeIndex_int) <= i_ch_cc;
            end if;
        end if;
      end process;

end Behavioral;
