library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity TuileBuffActor is
    Port(
    i_x : in STD_LOGIC_VECTOR (3 downto 0);
    i_y : in STD_LOGIC_VECTOR (3 downto 0);
    i_actor_is_present : in STD_LOGIC;
    i_tile_id : in STD_LOGIC_VECTOR (2 downto 0);
    i_ch_x : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_y : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_cc : in STD_LOGIC_VECTOR (3 downto 0);
    i_ch_we : in std_logic;
    i_clk : in STD_LOGIC;
    i_flip_y : in STD_LOGIC;
    i_tile_id_write : in STD_LOGIC_VECTOR (2 downto 0);
    o_is_actor_present : out std_logic;
    o_colorCode : out STD_LOGIC_VECTOR (3 downto 0));
end TuileBuffActor;

architecture Behavioral of TuileBuffActor is
constant wh : std_logic_vector (3 downto 0) := "0000"; -- White
constant bl : std_logic_vector (3 downto 0) := "0001"; -- Black
constant ye : std_logic_vector (3 downto 0) := "0010"; -- Yellow
constant dg : std_logic_vector (3 downto 0) := "0011"; -- Dark Green
constant oa : std_logic_vector (3 downto 0) := "0100"; -- Orange
constant bu : std_logic_vector (3 downto 0) := "0101"; -- Blue
constant ge : std_logic_vector (3 downto 0) := "0110"; -- Green
constant lo : std_logic_vector (3 downto 0) := "0111"; -- Light Brown
constant br : std_logic_vector (3 downto 0) := "1000"; -- Brown
constant lg : std_logic_vector (3 downto 0) := "1001"; -- Light Gray
constant gr : std_logic_vector (3 downto 0) := "1010"; -- Gray
constant lb : std_logic_vector (3 downto 0) := "1011"; -- Light Blue
constant sb : std_logic_vector (3 downto 0) := "1100"; -- Sky Blue
constant sa : std_logic_vector (3 downto 0) := "1101"; -- Salmon
constant pi : std_logic_vector (3 downto 0) := "1110"; -- Pink
constant pu : std_logic_vector (3 downto 0) := "1111"; -- darker green

    type tuile_out_array_t is array (0 to 7) of std_logic_vector(3 downto 0);
    signal tuile_outputs : tuile_out_array_t;
    signal tuile_write_enable : std_logic_vector(7 downto 0);
    
    type tile_d_array_t is array (0 to 2047) of std_logic_vector(3 downto 0);
    signal tile_data_map_d : tile_d_array_t :=
    (
0 => bl,
1 => bl,
2 => bl,
3 => bl,
4 => bl,
5 => pu,
6 => pu,
7 => pu,
8 => pu,
9 => pu,
10 => pu,
11 => pu,
12 => pu,
13 => pu,
14 => pu,
15 => pu,
16 => pu,
17 => pu,
18 => pu,
19 => pu,
20 => pu,
21 => pu,
22 => pu,
23 => bl,
24 => bl,
25 => bl,
26 => bl,
27 => bl,
28 => bl,
29 => bl,
30 => bl,
31 => bl,
32 => bl,
33 => bl,
34 => bl,
35 => bl,
36 => bl,
37 => bl,
38 => bl,
39 => bl,
40 => bl,
41 => bl,
42 => bl,
43 => bl,
44 => bl,
45 => bl,
46 => bl,
47 => bl,
48 => bl,
49 => bl,
50 => bl,
51 => bl,
52 => bl,
53 => bl,
54 => bl,
55 => bl,
56 => bl,
57 => bl,
58 => bl,
59 => bl,
60 => bl,
61 => bl,
62 => bl,
63 => bl,
64 => bl,
65 => bl,
66 => bl,
67 => bl,
68 => bl,
69 => bl,
70 => bl,
71 => bl,
72 => bl,
73 => bl,
74 => bl,
75 => bl,
76 => bl,
77 => bl,
78 => bl,
79 => bl,
80 => bl,
81 => bl,
82 => bl,
83 => bl,
84 => bl,
85 => bl,
86 => bl,
87 => bl,
88 => bl,
89 => bl,
90 => bl,
91 => bl,
92 => bl,
93 => bl,
94 => bl,
95 => bl,
96 => bl,
97 => bl,
98 => bl,
99 => bl,
100 => bl,
101 => bl,
102 => bl,
103 => bl,
104 => bl,
105 => bl,
106 => bl,
107 => bl,
108 => bl,
109 => bl,
110 => bl,
111 => bl,
112 => bl,
113 => bl,
114 => bl,
115 => bl,
116 => bl,
117 => bl,
118 => bl,
119 => bl,
120 => bl,
121 => bl,
122 => bl,
123 => bl,
124 => bl,
125 => bl,
126 => bl,
127 => bl,
128 => bl,
129 => bl,
130 => bl,
131 => bl,
132 => bl,
133 => bl,
134 => bl,
135 => bl,
136 => bl,
137 => bl,
138 => bl,
139 => bl,
140 => bl,
141 => bl,
142 => bl,
143 => bl,
144 => bl,
145 => bl,
146 => bl,
147 => bl,
148 => bl,
149 => bl,
150 => bl,
151 => bl,
152 => bl,
153 => bl,
154 => bl,
155 => bl,
156 => bl,
157 => bl,
158 => bl,
159 => bl,
160 => bl,
161 => bl,
162 => bl,
163 => bl,
164 => bl,
165 => bl,
166 => bl,
167 => bl,
168 => bl,
169 => bl,
170 => bl,
171 => bl,
172 => bl,
173 => bl,
174 => bl,
175 => bl,
176 => bl,
177 => bl,
178 => bl,
179 => bl,
180 => bl,
181 => bl,
182 => bl,
183 => bl,
184 => bl,
185 => bl,
186 => bl,
187 => bl,
188 => bl,
189 => bl,
190 => bl,
191 => bl,
192 => bl,
193 => bl,
194 => bl,
195 => bl,
196 => bl,
197 => bl,
198 => bl,
199 => bl,
200 => bl,
201 => bl,
202 => bl,
203 => bl,
204 => bl,
205 => bl,
206 => bl,
207 => bl,
208 => bl,
209 => bl,
210 => bl,
211 => bl,
212 => bl,
213 => bl,
214 => bl,
215 => bl,
216 => bl,
217 => bl,
218 => bl,
219 => bl,
220 => bl,
221 => bl,
222 => bl,
223 => bl,
224 => bl,
225 => bl,
226 => bl,
227 => bl,
228 => bl,
229 => bl,
230 => bl,
231 => bl,
232 => bl,
233 => bl,
234 => bl,
235 => bl,
236 => bl,
237 => bl,
238 => bl,
239 => bl,
240 => bl,
241 => bl,
242 => bl,
243 => bl,
244 => bl,
245 => bl,
246 => bl,
247 => bl,
248 => bl,
249 => bl,
250 => bl,
251 => bl,
252 => bl,
253 => bl,
254 => bl,
255 => bl,
256 => wh,
257 => wh,
258 => wh,
259 => wh,
260 => wh,
261 => wh,
262 => wh,
263 => wh,
264 => bu,
265 => wh,
266 => wh,
267 => wh,
268 => wh,
269 => wh,
270 => wh,
271 => wh,
272 => wh,
273 => wh,
274 => wh,
275 => wh,
276 => wh,
277 => wh,
278 => wh,
279 => bu,
280 => wh,
281 => wh,
282 => wh,
283 => wh,
284 => wh,
285 => wh,
286 => wh,
287 => wh,
288 => wh,
289 => wh,
290 => bl,
291 => wh,
292 => wh,
293 => wh,
294 => bu,
295 => wh,
296 => wh,
297 => wh,
298 => wh,
299 => wh,
300 => wh,
301 => wh,
302 => wh,
303 => wh,
304 => wh,
305 => bl,
306 => bl,
307 => bl,
308 => wh,
309 => bu,
310 => wh,
311 => wh,
312 => wh,
313 => wh,
314 => wh,
315 => wh,
316 => wh,
317 => wh,
318 => wh,
319 => wh,
320 => wh,
321 => bl,
322 => bl,
323 => bl,
324 => oa,
325 => wh,
326 => wh,
327 => wh,
328 => wh,
329 => wh,
330 => wh,
331 => wh,
332 => wh,
333 => wh,
334 => wh,
335 => wh,
336 => wh,
337 => wh,
338 => bl,
339 => oa,
340 => bl,
341 => wh,
342 => wh,
343 => wh,
344 => wh,
345 => wh,
346 => wh,
347 => wh,
348 => wh,
349 => wh,
350 => wh,
351 => wh,
352 => wh,
353 => wh,
354 => oa,
355 => bl,
356 => bl,
357 => bl,
358 => wh,
359 => wh,
360 => wh,
361 => wh,
362 => wh,
363 => wh,
364 => wh,
365 => wh,
366 => wh,
367 => wh,
368 => wh,
369 => bu,
370 => wh,
371 => bl,
372 => bl,
373 => bl,
374 => bl,
375 => wh,
376 => bl,
377 => bl,
378 => bl,
379 => bl,
380 => bl,
381 => bl,
382 => wh,
383 => bu,
384 => wh,
385 => bu,
386 => wh,
387 => wh,
388 => bl,
389 => bl,
390 => bl,
391 => bl,
392 => bl,
393 => bl,
394 => bl,
395 => bl,
396 => bl,
397 => bl,
398 => bu,
399 => wh,
400 => bu,
401 => wh,
402 => wh,
403 => wh,
404 => wh,
405 => bl,
406 => bl,
407 => bl,
408 => bl,
409 => bl,
410 => bl,
411 => bl,
412 => bl,
413 => bu,
414 => wh,
415 => wh,
416 => bu,
417 => wh,
418 => wh,
419 => wh,
420 => wh,
421 => wh,
422 => bl,
423 => bl,
424 => bl,
425 => bl,
426 => bl,
427 => bl,
428 => bu,
429 => wh,
430 => wh,
431 => wh,
432 => bu,
433 => wh,
434 => wh,
435 => wh,
436 => wh,
437 => wh,
438 => wh,
439 => bl,
440 => bl,
441 => bl,
442 => wh,
443 => bu,
444 => wh,
445 => wh,
446 => wh,
447 => wh,
448 => bu,
449 => wh,
450 => wh,
451 => wh,
452 => wh,
453 => wh,
454 => wh,
455 => wh,
456 => wh,
457 => wh,
458 => bu,
459 => wh,
460 => wh,
461 => wh,
462 => wh,
463 => wh,
464 => wh,
465 => bu,
466 => wh,
467 => wh,
468 => wh,
469 => wh,
470 => wh,
471 => wh,
472 => wh,
473 => bu,
474 => wh,
475 => wh,
476 => wh,
477 => wh,
478 => wh,
479 => wh,
480 => wh,
481 => wh,
482 => bu,
483 => wh,
484 => wh,
485 => wh,
486 => wh,
487 => bu,
488 => bu,
489 => wh,
490 => wh,
491 => wh,
492 => wh,
493 => wh,
494 => wh,
495 => wh,
496 => wh,
497 => wh,
498 => wh,
499 => bu,
500 => bu,
501 => bu,
502 => bu,
503 => wh,
504 => wh,
505 => wh,
506 => wh,
507 => wh,
508 => wh,
509 => wh,
510 => wh,
511 => wh,
512 => wh,
513 => wh,
514 => wh,
515 => wh,
516 => wh,
517 => wh,
518 => wh,
519 => wh,
520 => wh,
521 => bu,
522 => bu,
523 => bu,
524 => bu,
525 => wh,
526 => wh,
527 => bl,
528 => wh,
529 => wh,
530 => wh,
531 => wh,
532 => wh,
533 => wh,
534 => wh,
535 => bu,
536 => bu,
537 => wh,
538 => wh,
539 => wh,
540 => wh,
541 => bu,
542 => bl,
543 => bl,
544 => wh,
545 => wh,
546 => wh,
547 => wh,
548 => wh,
549 => wh,
550 => bu,
551 => wh,
552 => wh,
553 => wh,
554 => wh,
555 => wh,
556 => wh,
557 => oa,
558 => bl,
559 => bl,
560 => wh,
561 => wh,
562 => wh,
563 => wh,
564 => wh,
565 => bu,
566 => wh,
567 => wh,
568 => wh,
569 => wh,
570 => wh,
571 => wh,
572 => wh,
573 => bl,
574 => oa,
575 => bl,
576 => wh,
577 => wh,
578 => wh,
579 => wh,
580 => bu,
581 => wh,
582 => wh,
583 => wh,
584 => wh,
585 => wh,
586 => wh,
587 => wh,
588 => bl,
589 => bl,
590 => bl,
591 => bu,
592 => wh,
593 => wh,
594 => wh,
595 => bu,
596 => wh,
597 => wh,
598 => wh,
599 => wh,
600 => wh,
601 => wh,
602 => wh,
603 => bl,
604 => bl,
605 => bl,
606 => wh,
607 => bu,
608 => wh,
609 => wh,
610 => bu,
611 => wh,
612 => wh,
613 => wh,
614 => wh,
615 => wh,
616 => wh,
617 => bl,
618 => bl,
619 => bl,
620 => bl,
621 => bl,
622 => wh,
623 => bu,
624 => wh,
625 => bu,
626 => wh,
627 => wh,
628 => wh,
629 => wh,
630 => wh,
631 => bl,
632 => bl,
633 => bl,
634 => bl,
635 => bl,
636 => bl,
637 => wh,
638 => wh,
639 => bu,
640 => bu,
641 => wh,
642 => oa,
643 => oa,
644 => oa,
645 => oa,
646 => bl,
647 => bl,
648 => bl,
649 => bl,
650 => bl,
651 => bl,
652 => wh,
653 => wh,
654 => bu,
655 => wh,
656 => wh,
657 => oa,
658 => bl,
659 => bl,
660 => bl,
661 => bl,
662 => oa,
663 => bl,
664 => bl,
665 => bl,
666 => bl,
667 => wh,
668 => wh,
669 => bu,
670 => wh,
671 => wh,
672 => oa,
673 => bl,
674 => bl,
675 => bl,
676 => bl,
677 => bl,
678 => bl,
679 => oa,
680 => bl,
681 => bl,
682 => bl,
683 => wh,
684 => bu,
685 => wh,
686 => wh,
687 => wh,
688 => oa,
689 => bl,
690 => bl,
691 => bl,
692 => bl,
693 => bl,
694 => bl,
695 => oa,
696 => bl,
697 => bl,
698 => wh,
699 => bu,
700 => wh,
701 => wh,
702 => wh,
703 => wh,
704 => oa,
705 => bl,
706 => bl,
707 => bl,
708 => bl,
709 => bl,
710 => bl,
711 => oa,
712 => bl,
713 => wh,
714 => bu,
715 => wh,
716 => wh,
717 => wh,
718 => wh,
719 => wh,
720 => oa,
721 => bl,
722 => bl,
723 => bl,
724 => bl,
725 => bl,
726 => bl,
727 => oa,
728 => wh,
729 => bu,
730 => wh,
731 => wh,
732 => wh,
733 => wh,
734 => wh,
735 => wh,
736 => bl,
737 => oa,
738 => bl,
739 => bl,
740 => bl,
741 => bl,
742 => oa,
743 => wh,
744 => bu,
745 => wh,
746 => wh,
747 => wh,
748 => wh,
749 => wh,
750 => wh,
751 => wh,
752 => bl,
753 => bl,
754 => oa,
755 => oa,
756 => oa,
757 => oa,
758 => wh,
759 => bu,
760 => wh,
761 => wh,
762 => wh,
763 => wh,
764 => wh,
765 => wh,
766 => wh,
767 => wh,
768 => bl,
769 => bl,
770 => bl,
771 => bl,
772 => bl,
773 => bl,
774 => bl,
775 => bl,
776 => bl,
777 => bl,
778 => bl,
779 => bl,
780 => bl,
781 => bl,
782 => bl,
783 => bl,
784 => bl,
785 => bl,
786 => bl,
787 => bl,
788 => bl,
789 => bl,
790 => bl,
791 => bl,
792 => bl,
793 => bl,
794 => bl,
795 => bl,
796 => bl,
797 => bl,
798 => bl,
799 => bl,
800 => bl,
801 => bl,
802 => bl,
803 => bl,
804 => bl,
805 => bl,
806 => bl,
807 => bl,
808 => bl,
809 => bl,
810 => bl,
811 => bl,
812 => bl,
813 => bl,
814 => bl,
815 => bl,
816 => bl,
817 => bl,
818 => bl,
819 => bl,
820 => bl,
821 => bl,
822 => bl,
823 => bl,
824 => bl,
825 => bl,
826 => bl,
827 => bl,
828 => bl,
829 => bl,
830 => bl,
831 => bl,
832 => bl,
833 => bl,
834 => bl,
835 => bl,
836 => bl,
837 => bl,
838 => bl,
839 => bl,
840 => bl,
841 => bl,
842 => bl,
843 => bl,
844 => bl,
845 => bl,
846 => bl,
847 => bl,
848 => bl,
849 => bl,
850 => bl,
851 => bl,
852 => bl,
853 => bl,
854 => bl,
855 => bl,
856 => bl,
857 => bl,
858 => bl,
859 => bl,
860 => bl,
861 => bl,
862 => bl,
863 => bl,
864 => bl,
865 => bl,
866 => bl,
867 => bl,
868 => bl,
869 => bl,
870 => bl,
871 => bl,
872 => bl,
873 => bl,
874 => bl,
875 => bl,
876 => bl,
877 => bl,
878 => bl,
879 => bl,
880 => bl,
881 => bl,
882 => bl,
883 => bl,
884 => bl,
885 => bl,
886 => bl,
887 => bl,
888 => bl,
889 => bl,
890 => bl,
891 => bl,
892 => bl,
893 => bl,
894 => bl,
895 => bl,
896 => bl,
897 => bl,
898 => bl,
899 => bl,
900 => bl,
901 => bl,
902 => bl,
903 => bl,
904 => bl,
905 => bl,
906 => bl,
907 => bl,
908 => bl,
909 => bl,
910 => bl,
911 => bl,
912 => bl,
913 => bl,
914 => bl,
915 => bl,
916 => bl,
917 => bl,
918 => bl,
919 => bl,
920 => bl,
921 => bl,
922 => bl,
923 => bl,
924 => bl,
925 => bl,
926 => bl,
927 => bl,
928 => bl,
929 => bl,
930 => bl,
931 => bl,
932 => bl,
933 => bl,
934 => bl,
935 => bl,
936 => bl,
937 => bl,
938 => bl,
939 => bl,
940 => bl,
941 => bl,
942 => bl,
943 => bl,
944 => bl,
945 => bl,
946 => bl,
947 => bl,
948 => bl,
949 => bl,
950 => bl,
951 => bl,
952 => bl,
953 => bl,
954 => bl,
955 => bl,
956 => bl,
957 => bl,
958 => bl,
959 => bl,
960 => bl,
961 => bl,
962 => bl,
963 => bl,
964 => bl,
965 => bl,
966 => bl,
967 => bl,
968 => bl,
969 => bl,
970 => bl,
971 => bl,
972 => bl,
973 => bl,
974 => bl,
975 => bl,
976 => bl,
977 => bl,
978 => bl,
979 => bl,
980 => bl,
981 => bl,
982 => bl,
983 => bl,
984 => bl,
985 => bl,
986 => bl,
987 => bl,
988 => bl,
989 => bl,
990 => bl,
991 => bl,
992 => bl,
993 => bl,
994 => bl,
995 => bl,
996 => bl,
997 => bl,
998 => bl,
999 => bl,
1000 => bl,
1001 => bl,
1002 => bl,
1003 => bl,
1004 => bl,
1005 => bl,
1006 => bl,
1007 => bl,
1008 => bl,
1009 => bl,
1010 => bl,
1011 => bl,
1012 => bl,
1013 => bl,
1014 => bl,
1015 => bl,
1016 => bl,
1017 => bl,
1018 => bl,
1019 => bl,
1020 => bl,
1021 => bl,
1022 => bl,
1023 => bl,
1024 => bl,
1025 => bl,
1026 => bl,
1027 => bl,
1028 => bl,
1029 => bl,
1030 => bl,
1031 => bl,
1032 => bl,
1033 => bl,
1034 => bl,
1035 => bl,
1036 => bl,
1037 => bl,
1038 => bl,
1039 => bl,
1040 => bl,
1041 => bl,
1042 => bl,
1043 => bl,
1044 => bl,
1045 => bl,
1046 => bl,
1047 => bl,
1048 => bl,
1049 => bl,
1050 => bl,
1051 => bl,
1052 => bl,
1053 => bl,
1054 => bl,
1055 => bl,
1056 => bl,
1057 => bl,
1058 => bl,
1059 => bl,
1060 => bl,
1061 => bl,
1062 => bl,
1063 => bl,
1064 => bl,
1065 => bl,
1066 => bl,
1067 => bl,
1068 => bl,
1069 => bl,
1070 => bl,
1071 => bl,
1072 => bl,
1073 => bl,
1074 => bl,
1075 => bl,
1076 => bl,
1077 => bl,
1078 => bl,
1079 => bl,
1080 => bl,
1081 => bl,
1082 => bl,
1083 => bl,
1084 => bl,
1085 => bl,
1086 => bl,
1087 => bl,
1088 => bl,
1089 => bl,
1090 => bl,
1091 => bl,
1092 => bl,
1093 => bl,
1094 => bl,
1095 => bl,
1096 => bl,
1097 => bl,
1098 => bl,
1099 => bl,
1100 => bl,
1101 => bl,
1102 => bl,
1103 => bl,
1104 => bl,
1105 => bl,
1106 => bl,
1107 => bl,
1108 => bl,
1109 => bl,
1110 => bl,
1111 => bl,
1112 => bl,
1113 => bl,
1114 => bl,
1115 => bl,
1116 => bl,
1117 => bl,
1118 => bl,
1119 => bl,
1120 => bl,
1121 => bl,
1122 => bl,
1123 => bl,
1124 => bl,
1125 => bl,
1126 => bl,
1127 => bl,
1128 => bl,
1129 => bl,
1130 => bl,
1131 => bl,
1132 => bl,
1133 => bl,
1134 => bl,
1135 => bl,
1136 => bl,
1137 => bl,
1138 => bl,
1139 => bl,
1140 => bl,
1141 => bl,
1142 => bl,
1143 => bl,
1144 => bl,
1145 => bl,
1146 => bl,
1147 => bl,
1148 => bl,
1149 => bl,
1150 => bl,
1151 => bl,
1152 => bl,
1153 => bl,
1154 => bl,
1155 => bl,
1156 => bl,
1157 => bl,
1158 => bl,
1159 => bl,
1160 => bl,
1161 => bl,
1162 => bl,
1163 => bl,
1164 => bl,
1165 => bl,
1166 => bl,
1167 => bl,
1168 => bl,
1169 => bl,
1170 => bl,
1171 => bl,
1172 => bl,
1173 => bl,
1174 => bl,
1175 => bl,
1176 => bl,
1177 => bl,
1178 => bl,
1179 => bl,
1180 => bl,
1181 => bl,
1182 => bl,
1183 => bl,
1184 => bl,
1185 => bl,
1186 => bl,
1187 => bl,
1188 => bl,
1189 => bl,
1190 => bl,
1191 => bl,
1192 => bl,
1193 => bl,
1194 => bl,
1195 => bl,
1196 => bl,
1197 => bl,
1198 => bl,
1199 => bl,
1200 => bl,
1201 => bl,
1202 => bl,
1203 => bl,
1204 => bl,
1205 => bl,
1206 => bl,
1207 => bl,
1208 => bl,
1209 => bl,
1210 => bl,
1211 => bl,
1212 => bl,
1213 => bl,
1214 => bl,
1215 => bl,
1216 => bl,
1217 => bl,
1218 => bl,
1219 => bl,
1220 => bl,
1221 => bl,
1222 => bl,
1223 => bl,
1224 => bl,
1225 => bl,
1226 => bl,
1227 => bl,
1228 => bl,
1229 => bl,
1230 => bl,
1231 => bl,
1232 => bl,
1233 => bl,
1234 => bl,
1235 => bl,
1236 => bl,
1237 => bl,
1238 => bl,
1239 => bl,
1240 => bl,
1241 => bl,
1242 => bl,
1243 => bl,
1244 => bl,
1245 => bl,
1246 => bl,
1247 => bl,
1248 => bl,
1249 => bl,
1250 => bl,
1251 => bl,
1252 => bl,
1253 => bl,
1254 => bl,
1255 => bl,
1256 => bl,
1257 => bl,
1258 => bl,
1259 => bl,
1260 => bl,
1261 => bl,
1262 => bl,
1263 => bl,
1264 => bl,
1265 => bl,
1266 => bl,
1267 => bl,
1268 => bl,
1269 => bl,
1270 => bl,
1271 => bl,
1272 => bl,
1273 => bl,
1274 => bl,
1275 => bl,
1276 => bl,
1277 => bl,
1278 => bl,
1279 => bl,
1280 => bl,
1281 => bl,
1282 => bl,
1283 => bl,
1284 => bl,
1285 => bl,
1286 => bl,
1287 => bl,
1288 => bl,
1289 => bl,
1290 => bl,
1291 => bl,
1292 => bl,
1293 => bl,
1294 => bl,
1295 => bl,
1296 => bl,
1297 => bl,
1298 => bl,
1299 => bl,
1300 => bl,
1301 => bl,
1302 => bl,
1303 => bl,
1304 => bl,
1305 => bl,
1306 => bl,
1307 => bl,
1308 => bl,
1309 => bl,
1310 => bl,
1311 => bl,
1312 => bl,
1313 => bl,
1314 => bl,
1315 => bl,
1316 => bl,
1317 => bl,
1318 => bl,
1319 => bl,
1320 => bl,
1321 => bl,
1322 => bl,
1323 => bl,
1324 => bl,
1325 => bl,
1326 => bl,
1327 => bl,
1328 => bl,
1329 => bl,
1330 => bl,
1331 => bl,
1332 => bl,
1333 => bl,
1334 => bl,
1335 => bl,
1336 => bl,
1337 => bl,
1338 => bl,
1339 => bl,
1340 => bl,
1341 => bl,
1342 => bl,
1343 => bl,
1344 => bl,
1345 => bl,
1346 => bl,
1347 => bl,
1348 => bl,
1349 => bl,
1350 => bl,
1351 => bl,
1352 => bl,
1353 => bl,
1354 => bl,
1355 => bl,
1356 => bl,
1357 => bl,
1358 => bl,
1359 => bl,
1360 => bl,
1361 => bl,
1362 => bl,
1363 => bl,
1364 => bl,
1365 => bl,
1366 => bl,
1367 => bl,
1368 => bl,
1369 => bl,
1370 => bl,
1371 => bl,
1372 => bl,
1373 => bl,
1374 => bl,
1375 => bl,
1376 => bl,
1377 => bl,
1378 => bl,
1379 => bl,
1380 => bl,
1381 => bl,
1382 => bl,
1383 => bl,
1384 => bl,
1385 => bl,
1386 => bl,
1387 => bl,
1388 => bl,
1389 => bl,
1390 => bl,
1391 => bl,
1392 => bl,
1393 => bl,
1394 => bl,
1395 => bl,
1396 => bl,
1397 => bl,
1398 => bl,
1399 => bl,
1400 => bl,
1401 => bl,
1402 => bl,
1403 => bl,
1404 => bl,
1405 => bl,
1406 => bl,
1407 => bl,
1408 => bl,
1409 => bl,
1410 => bl,
1411 => bl,
1412 => bl,
1413 => bl,
1414 => bl,
1415 => bl,
1416 => bl,
1417 => bl,
1418 => bl,
1419 => bl,
1420 => bl,
1421 => bl,
1422 => bl,
1423 => bl,
1424 => bl,
1425 => bl,
1426 => bl,
1427 => bl,
1428 => bl,
1429 => bl,
1430 => bl,
1431 => bl,
1432 => bl,
1433 => bl,
1434 => bl,
1435 => bl,
1436 => bl,
1437 => bl,
1438 => bl,
1439 => bl,
1440 => bl,
1441 => bl,
1442 => bl,
1443 => bl,
1444 => bl,
1445 => bl,
1446 => bl,
1447 => bl,
1448 => bl,
1449 => bl,
1450 => bl,
1451 => bl,
1452 => bl,
1453 => bl,
1454 => bl,
1455 => bl,
1456 => bl,
1457 => bl,
1458 => bl,
1459 => bl,
1460 => bl,
1461 => bl,
1462 => bl,
1463 => bl,
1464 => bl,
1465 => bl,
1466 => bl,
1467 => bl,
1468 => bl,
1469 => bl,
1470 => bl,
1471 => bl,
1472 => bl,
1473 => bl,
1474 => bl,
1475 => bl,
1476 => bl,
1477 => bl,
1478 => bl,
1479 => bl,
1480 => bl,
1481 => bl,
1482 => bl,
1483 => bl,
1484 => bl,
1485 => bl,
1486 => bl,
1487 => bl,
1488 => bl,
1489 => bl,
1490 => bl,
1491 => bl,
1492 => bl,
1493 => bl,
1494 => bl,
1495 => bl,
1496 => bl,
1497 => bl,
1498 => bl,
1499 => bl,
1500 => bl,
1501 => bl,
1502 => bl,
1503 => bl,
1504 => bl,
1505 => bl,
1506 => bl,
1507 => bl,
1508 => bl,
1509 => bl,
1510 => bl,
1511 => bl,
1512 => bl,
1513 => bl,
1514 => bl,
1515 => bl,
1516 => bl,
1517 => bl,
1518 => bl,
1519 => bl,
1520 => bl,
1521 => bl,
1522 => bl,
1523 => bl,
1524 => bl,
1525 => bl,
1526 => bl,
1527 => bl,
1528 => bl,
1529 => bl,
1530 => bl,
1531 => bl,
1532 => bl,
1533 => bl,
1534 => bl,
1535 => bl,
1536 => bl,
1537 => bl,
1538 => bl,
1539 => bl,
1540 => bl,
1541 => bl,
1542 => bl,
1543 => bl,
1544 => bl,
1545 => bl,
1546 => bl,
1547 => bl,
1548 => bl,
1549 => bl,
1550 => bl,
1551 => bl,
1552 => bl,
1553 => bl,
1554 => bl,
1555 => bl,
1556 => bl,
1557 => bl,
1558 => bl,
1559 => bl,
1560 => bl,
1561 => bl,
1562 => bl,
1563 => bl,
1564 => bl,
1565 => bl,
1566 => bl,
1567 => bl,
1568 => bl,
1569 => bl,
1570 => bl,
1571 => bl,
1572 => bl,
1573 => bl,
1574 => bl,
1575 => bl,
1576 => bl,
1577 => bl,
1578 => bl,
1579 => bl,
1580 => bl,
1581 => bl,
1582 => bl,
1583 => bl,
1584 => bl,
1585 => bl,
1586 => bl,
1587 => bl,
1588 => bl,
1589 => bl,
1590 => bl,
1591 => bl,
1592 => bl,
1593 => bl,
1594 => bl,
1595 => bl,
1596 => bl,
1597 => bl,
1598 => bl,
1599 => bl,
1600 => bl,
1601 => bl,
1602 => bl,
1603 => bl,
1604 => bl,
1605 => bl,
1606 => bl,
1607 => bl,
1608 => bl,
1609 => bl,
1610 => bl,
1611 => bl,
1612 => bl,
1613 => bl,
1614 => bl,
1615 => bl,
1616 => bl,
1617 => bl,
1618 => bl,
1619 => bl,
1620 => bl,
1621 => bl,
1622 => bl,
1623 => bl,
1624 => bl,
1625 => bl,
1626 => bl,
1627 => bl,
1628 => bl,
1629 => bl,
1630 => bl,
1631 => bl,
1632 => bl,
1633 => bl,
1634 => bl,
1635 => bl,
1636 => bl,
1637 => bl,
1638 => bl,
1639 => bl,
1640 => bl,
1641 => bl,
1642 => bl,
1643 => bl,
1644 => bl,
1645 => bl,
1646 => bl,
1647 => bl,
1648 => bl,
1649 => bl,
1650 => bl,
1651 => bl,
1652 => bl,
1653 => bl,
1654 => bl,
1655 => bl,
1656 => bl,
1657 => bl,
1658 => bl,
1659 => bl,
1660 => bl,
1661 => bl,
1662 => bl,
1663 => bl,
1664 => bl,
1665 => bl,
1666 => bl,
1667 => bl,
1668 => bl,
1669 => bl,
1670 => bl,
1671 => bl,
1672 => bl,
1673 => bl,
1674 => bl,
1675 => bl,
1676 => bl,
1677 => bl,
1678 => bl,
1679 => bl,
1680 => bl,
1681 => bl,
1682 => bl,
1683 => bl,
1684 => bl,
1685 => bl,
1686 => bl,
1687 => bl,
1688 => bl,
1689 => bl,
1690 => bl,
1691 => bl,
1692 => bl,
1693 => bl,
1694 => bl,
1695 => bl,
1696 => bl,
1697 => bl,
1698 => bl,
1699 => bl,
1700 => bl,
1701 => bl,
1702 => bl,
1703 => bl,
1704 => bl,
1705 => bl,
1706 => bl,
1707 => bl,
1708 => bl,
1709 => bl,
1710 => bl,
1711 => bl,
1712 => bl,
1713 => bl,
1714 => bl,
1715 => bl,
1716 => bl,
1717 => bl,
1718 => bl,
1719 => bl,
1720 => bl,
1721 => bl,
1722 => bl,
1723 => bl,
1724 => bl,
1725 => bl,
1726 => bl,
1727 => bl,
1728 => bl,
1729 => bl,
1730 => bl,
1731 => bl,
1732 => bl,
1733 => bl,
1734 => bl,
1735 => bl,
1736 => bl,
1737 => bl,
1738 => bl,
1739 => bl,
1740 => bl,
1741 => bl,
1742 => bl,
1743 => bl,
1744 => bl,
1745 => bl,
1746 => bl,
1747 => bl,
1748 => bl,
1749 => bl,
1750 => bl,
1751 => bl,
1752 => bl,
1753 => bl,
1754 => bl,
1755 => bl,
1756 => bl,
1757 => bl,
1758 => bl,
1759 => bl,
1760 => bl,
1761 => bl,
1762 => bl,
1763 => bl,
1764 => bl,
1765 => bl,
1766 => bl,
1767 => bl,
1768 => bl,
1769 => bl,
1770 => bl,
1771 => bl,
1772 => bl,
1773 => bl,
1774 => bl,
1775 => bl,
1776 => bl,
1777 => bl,
1778 => bl,
1779 => bl,
1780 => bl,
1781 => bl,
1782 => bl,
1783 => bl,
1784 => bl,
1785 => bl,
1786 => bl,
1787 => bl,
1788 => bl,
1789 => bl,
1790 => bl,
1791 => bl,
1792 => bl,
1793 => bl,
1794 => bl,
1795 => bl,
1796 => bl,
1797 => bl,
1798 => bl,
1799 => bl,
1800 => bl,
1801 => bl,
1802 => bl,
1803 => bl,
1804 => bl,
1805 => bl,
1806 => bl,
1807 => bl,
1808 => bl,
1809 => bl,
1810 => bl,
1811 => bl,
1812 => bl,
1813 => bl,
1814 => bl,
1815 => bl,
1816 => bl,
1817 => bl,
1818 => bl,
1819 => bl,
1820 => bl,
1821 => bl,
1822 => bl,
1823 => bl,
1824 => bl,
1825 => bl,
1826 => bl,
1827 => bl,
1828 => bl,
1829 => bl,
1830 => bl,
1831 => bl,
1832 => bl,
1833 => bl,
1834 => bl,
1835 => bl,
1836 => bl,
1837 => bl,
1838 => bl,
1839 => bl,
1840 => bl,
1841 => bl,
1842 => bl,
1843 => bl,
1844 => bl,
1845 => bl,
1846 => bl,
1847 => bl,
1848 => bl,
1849 => bl,
1850 => bl,
1851 => bl,
1852 => bl,
1853 => bl,
1854 => bl,
1855 => bl,
1856 => bl,
1857 => bl,
1858 => bl,
1859 => bl,
1860 => bl,
1861 => bl,
1862 => bl,
1863 => bl,
1864 => bl,
1865 => bl,
1866 => bl,
1867 => bl,
1868 => bl,
1869 => bl,
1870 => bl,
1871 => bl,
1872 => bl,
1873 => bl,
1874 => bl,
1875 => bl,
1876 => bl,
1877 => bl,
1878 => bl,
1879 => bl,
1880 => bl,
1881 => bl,
1882 => bl,
1883 => bl,
1884 => bl,
1885 => bl,
1886 => bl,
1887 => bl,
1888 => bl,
1889 => bl,
1890 => bl,
1891 => bl,
1892 => bl,
1893 => bl,
1894 => bl,
1895 => bl,
1896 => bl,
1897 => bl,
1898 => bl,
1899 => bl,
1900 => bl,
1901 => bl,
1902 => bl,
1903 => bl,
1904 => bl,
1905 => bl,
1906 => bl,
1907 => bl,
1908 => bl,
1909 => bl,
1910 => bl,
1911 => bl,
1912 => bl,
1913 => bl,
1914 => bl,
1915 => bl,
1916 => bl,
1917 => bl,
1918 => bl,
1919 => bl,
1920 => bl,
1921 => bl,
1922 => bl,
1923 => bl,
1924 => bl,
1925 => bl,
1926 => bl,
1927 => bl,
1928 => bl,
1929 => bl,
1930 => bl,
1931 => bl,
1932 => bl,
1933 => bl,
1934 => bl,
1935 => bl,
1936 => bl,
1937 => bl,
1938 => bl,
1939 => bl,
1940 => bl,
1941 => bl,
1942 => bl,
1943 => bl,
1944 => bl,
1945 => bl,
1946 => bl,
1947 => bl,
1948 => bl,
1949 => bl,
1950 => bl,
1951 => bl,
1952 => bl,
1953 => bl,
1954 => bl,
1955 => bl,
1956 => bl,
1957 => bl,
1958 => bl,
1959 => bl,
1960 => bl,
1961 => bl,
1962 => bl,
1963 => bl,
1964 => bl,
1965 => bl,
1966 => bl,
1967 => bl,
1968 => bl,
1969 => bl,
1970 => bl,
1971 => bl,
1972 => bl,
1973 => bl,
1974 => bl,
1975 => bl,
1976 => bl,
1977 => bl,
1978 => bl,
1979 => bl,
1980 => bl,
1981 => bl,
1982 => bl,
1983 => bl,
1984 => bl,
1985 => bl,
1986 => bl,
1987 => bl,
1988 => bl,
1989 => bl,
1990 => bl,
1991 => bl,
1992 => bl,
1993 => bl,
1994 => bl,
1995 => bl,
1996 => bl,
1997 => bl,
1998 => bl,
1999 => bl,
2000 => bl,
2001 => bl,
2002 => bl,
2003 => bl,
2004 => bl,
2005 => bl,
2006 => bl,
2007 => bl,
2008 => bl,
2009 => bl,
2010 => bl,
2011 => bl,
2012 => bl,
2013 => bl,
2014 => bl,
2015 => bl,
2016 => bl,
2017 => bl,
2018 => bl,
2019 => bl,
2020 => bl,
2021 => bl,
2022 => bl,
2023 => bl,
2024 => bl,
2025 => bl,
2026 => bl,
2027 => bl,
2028 => bl,
2029 => bl,
2030 => bl,
2031 => bl,
2032 => bl,
2033 => bl,
2034 => bl,
2035 => bl,
2036 => bl,
2037 => bl,
2038 => bl,
2039 => bl,
2040 => bl,
2041 => bl,
2042 => bl,
2043 => bl,
2044 => bl,
2045 => bl,
2046 => bl,
2047 => bl
    ); 
    
    attribute ram_style : string;
    attribute ram_style of tile_data_map_d : signal is "block";
begin
    
      process(i_tile_id, i_x, i_y)
          variable readIndex : std_logic_vector (10 downto 0);
          variable readIndex_int : integer;
          variable transparent : std_logic;
          variable readTuile : std_logic_vector (3 downto 0);
          begin
          readIndex := i_tile_id & i_y & i_x;
          readIndex_int := to_integer(unsigned(readIndex));
          readTuile := tile_data_map_d(readIndex_int);
          if readTuile = pu then
            o_is_actor_present <= '0';
          elsif i_actor_is_present = '1' then
            o_is_actor_present <= '1';
          end if;
          o_colorCode <= readTuile;
      end process;
      
      process(i_clk)
      variable writeIndex : std_logic_vector (10 downto 0);
      variable writeIndex_int : integer;
      begin
        if rising_edge(i_clk) then
            if i_ch_we = '1' then
                writeIndex := i_tile_id_write & i_ch_y & i_ch_x;
                writeIndex_int := to_integer(unsigned(writeIndex));
                tile_data_map_d(writeIndex_int) <= i_ch_cc;
            end if;
        end if;
      end process;

end Behavioral;
